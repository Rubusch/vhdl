// demo_diagnostic.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module demo_diagnostic (
		output wire [7:0] button_pio_export,    //    button_pio.export
		input  wire       clk_clk,              //           clk.clk
		output wire       lcd_display_RS,       //   lcd_display.RS
		output wire       lcd_display_RW,       //              .RW
		inout  wire [7:0] lcd_display_data,     //              .data
		output wire       lcd_display_E,        //              .E
		output wire [7:0] led_pio_export,       //       led_pio.export
		output wire [7:0] seven_seg_pio_export  // seven_seg_pio.export
	);

	wire         nios2_debug_reset_request_reset;                           // nios2:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                             // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [19:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [19:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_readdata;      // lcd_16207_0:readdata -> mm_interconnect_0:lcd_16207_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_16207_0_control_slave_address;       // mm_interconnect_0:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_0_lcd_16207_0_control_slave_read;          // mm_interconnect_0:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire         mm_interconnect_0_lcd_16207_0_control_slave_begintransfer; // mm_interconnect_0:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_0_lcd_16207_0_control_slave_write;         // mm_interconnect_0:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_writedata;     // mm_interconnect_0:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;          // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;       // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;           // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;              // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;             // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                         // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                       // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [2:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_seven_seg_s1_chipselect;                 // mm_interconnect_0:seven_seg_s1_chipselect -> seven_seg:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_s1_readdata;                   // seven_seg:readdata -> mm_interconnect_0:seven_seg_s1_readdata
	wire   [2:0] mm_interconnect_0_seven_seg_s1_address;                    // mm_interconnect_0:seven_seg_s1_address -> seven_seg:address
	wire         mm_interconnect_0_seven_seg_s1_write;                      // mm_interconnect_0:seven_seg_s1_write -> seven_seg:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_s1_writedata;                  // mm_interconnect_0:seven_seg_s1_writedata -> seven_seg:writedata
	wire         mm_interconnect_0_button_s1_chipselect;                    // mm_interconnect_0:button_s1_chipselect -> button:chipselect
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                      // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [2:0] mm_interconnect_0_button_s1_address;                       // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_button_s1_write;                         // mm_interconnect_0:button_s1_write -> button:write_n
	wire  [31:0] mm_interconnect_0_button_s1_writedata;                     // mm_interconnect_0:button_s1_writedata -> button:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_irq_irq;                                             // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [button:reset_n, irq_mapper:reset, jtag_uart:rst_n, lcd_16207_0:reset_n, led:reset_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, ram:reset, rst_translator:in_reset, seven_seg:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2:reset_req, ram:reset_req, rst_translator:reset_req_in]

	demo_diagnostic_button button (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.out_port   (button_pio_export)                       // external_connection.export
	);

	demo_diagnostic_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	demo_diagnostic_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (clk_clk),                                                   //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_display_RS),                                            //      external.export
		.LCD_RW        (lcd_display_RW),                                            //              .export
		.LCD_data      (lcd_display_data),                                          //              .export
		.LCD_E         (lcd_display_E)                                              //              .export
	);

	demo_diagnostic_button led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                       // external_connection.export
	);

	demo_diagnostic_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	demo_diagnostic_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	demo_diagnostic_button seven_seg (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_pio_export)                       // external_connection.export
	);

	demo_diagnostic_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                           clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address               (nios2_data_master_address),                                 //                 nios2_data_master.address
		.nios2_data_master_waitrequest           (nios2_data_master_waitrequest),                             //                                  .waitrequest
		.nios2_data_master_byteenable            (nios2_data_master_byteenable),                              //                                  .byteenable
		.nios2_data_master_read                  (nios2_data_master_read),                                    //                                  .read
		.nios2_data_master_readdata              (nios2_data_master_readdata),                                //                                  .readdata
		.nios2_data_master_write                 (nios2_data_master_write),                                   //                                  .write
		.nios2_data_master_writedata             (nios2_data_master_writedata),                               //                                  .writedata
		.nios2_data_master_debugaccess           (nios2_data_master_debugaccess),                             //                                  .debugaccess
		.nios2_instruction_master_address        (nios2_instruction_master_address),                          //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                      //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),                             //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),                         //                                  .readdata
		.button_s1_address                       (mm_interconnect_0_button_s1_address),                       //                         button_s1.address
		.button_s1_write                         (mm_interconnect_0_button_s1_write),                         //                                  .write
		.button_s1_readdata                      (mm_interconnect_0_button_s1_readdata),                      //                                  .readdata
		.button_s1_writedata                     (mm_interconnect_0_button_s1_writedata),                     //                                  .writedata
		.button_s1_chipselect                    (mm_interconnect_0_button_s1_chipselect),                    //                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.lcd_16207_0_control_slave_address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //         lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //                                  .write
		.lcd_16207_0_control_slave_read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //                                  .read
		.lcd_16207_0_control_slave_readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //                                  .readdata
		.lcd_16207_0_control_slave_writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //                                  .writedata
		.lcd_16207_0_control_slave_begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), //                                  .begintransfer
		.led_s1_address                          (mm_interconnect_0_led_s1_address),                          //                            led_s1.address
		.led_s1_write                            (mm_interconnect_0_led_s1_write),                            //                                  .write
		.led_s1_readdata                         (mm_interconnect_0_led_s1_readdata),                         //                                  .readdata
		.led_s1_writedata                        (mm_interconnect_0_led_s1_writedata),                        //                                  .writedata
		.led_s1_chipselect                       (mm_interconnect_0_led_s1_chipselect),                       //                                  .chipselect
		.nios2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),           //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),             //                                  .write
		.nios2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),              //                                  .read
		.nios2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),          //                                  .readdata
		.nios2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),         //                                  .writedata
		.nios2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),        //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),       //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),       //                                  .debugaccess
		.ram_s1_address                          (mm_interconnect_0_ram_s1_address),                          //                            ram_s1.address
		.ram_s1_write                            (mm_interconnect_0_ram_s1_write),                            //                                  .write
		.ram_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                         //                                  .readdata
		.ram_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                        //                                  .writedata
		.ram_s1_byteenable                       (mm_interconnect_0_ram_s1_byteenable),                       //                                  .byteenable
		.ram_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                       //                                  .chipselect
		.ram_s1_clken                            (mm_interconnect_0_ram_s1_clken),                            //                                  .clken
		.seven_seg_s1_address                    (mm_interconnect_0_seven_seg_s1_address),                    //                      seven_seg_s1.address
		.seven_seg_s1_write                      (mm_interconnect_0_seven_seg_s1_write),                      //                                  .write
		.seven_seg_s1_readdata                   (mm_interconnect_0_seven_seg_s1_readdata),                   //                                  .readdata
		.seven_seg_s1_writedata                  (mm_interconnect_0_seven_seg_s1_writedata),                  //                                  .writedata
		.seven_seg_s1_chipselect                 (mm_interconnect_0_seven_seg_s1_chipselect)                  //                                  .chipselect
	);

	demo_diagnostic_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_debug_reset_request_reset),    // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
