--
--  A[3..0] +-------+
--  --------| TWO   | C[3..0]
--  B[3..0] | INPUT |-------->
--  --------| MUXER |
--          +-------+
--              A
--              |
--  SEL --------+
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY QUADMUX IS
PORT( A   : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      B   : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      SEL : IN STD_LOGIC;
      C   : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) );
END ENTITY QUADMUX;


ARCHITECTURE QUADMUX_ARCH OF QUADMUX IS
BEGIN
-- A FIRST APPROACH (WORKING)
--	C <= A WHEN SEL = '0' ELSE B;

-- SYNTACTICALLY MORE ELEGANT TO USE SELECT IN CONTEXT OF A MULTIPLEXER
  WITH SEL SELECT
    C <= A WHEN '0',
         B WHEN OTHERS;
END ARCHITECTURE QUADMUX_ARCH;
