--
--
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SHIFTER_ENT IS
PORT( D : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
	; C : IN STD_LOGIC
	; S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END ENTITY SHIFTER_ENT;

ARCHITECTURE SHIFTER_ARCH OF SHIFTER_ENT IS
BEGIN

END ARCHITECTURE SHIFTER_ARCH;