-- hw adaptation for DE1SoC Board: fsm
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_FSM IS
PORT( CLK50 : IN STD_LOGIC
    ; KEY : IN STD_LOGIC
    ; SW  : IN STD_LOGIC_VECTOR(2 DOWNTO 0)
    ; LED : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END DE1SOC_FSM;

ARCHITECTURE DE1SOC OF DE1SOC_FSM IS
    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';
    SIGNAL KEYS : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
    SIGNAL LEDS : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');

BEGIN

    FSM_UNIT : ENTITY WORK.FSM
        PORT MAP(CLK => CLK, RST => RST, KEY => KEYS, LED => LEDS);

    -- IN
    CLK <= CLK50;
    RST <= NOT KEY;
    KEYS <= SW;

    -- OUT
    LED <= LEDS;

END DE1SOC;

