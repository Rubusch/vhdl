-- tb: alu
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_ALU IS
END TB_ALU;

ARCHITECTURE TB OF TB_ALU IS
    SIGNAL INVA : STD_LOGIC := '0';
    SIGNAL A : STD_LOGIC := '0';
    SIGNAL ENA : STD_LOGIC := '0';
    SIGNAL B : STD_LOGIC := '0';
    SIGNAL ENB : STD_LOGIC := '0';
    SIGNAL F : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL CARRY_IN : STD_LOGIC := '0';
    SIGNAL CARRY_OUT : STD_LOGIC := '0';
    SIGNAL CARRY_OUT_EXPECT : STD_LOGIC := '0';
    SIGNAL OUTPUT : STD_LOGIC := '0';
    SIGNAL OUTPUT_EXPECT : STD_LOGIC := '0';
    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    ALU_UNIT : ENTITY WORK.ALU
        PORT MAP (INVA => INVA
            , A => A
            , ENA => ENA
            , B => B
            , ENB => ENB
            , F => F
            , CARRY_IN => CARRY_IN
            , CARRY_OUT => CARRY_OUT
            , OUTPUT => OUTPUT
        );

    PROCESS
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE GOOD_NUM : BOOLEAN;
        VARIABLE SEPARATOR : CHARACTER;
        VARIABLE INPUT_INVA : STD_LOGIC;
        VARIABLE INPUT_A : STD_LOGIC;
        VARIABLE INPUT_ENA : STD_LOGIC;
        VARIABLE INPUT_B : STD_LOGIC;
        VARIABLE INPUT_ENB : STD_LOGIC;
        VARIABLE INPUT_F : STD_LOGIC_VECTOR(1 DOWNTO 0);
        VARIABLE INPUT_CARRY_IN : STD_LOGIC;
        VARIABLE INPUT_CARRY_OUT : STD_LOGIC;
        VARIABLE INPUT_OUTPUT : STD_LOGIC;
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("INVA,A,ENA,B,ENB,F,CARRY_IN,CARRY_OUT,CARRY_OUT_EXPECT,OUTPUT,OUTPUT_EXPECT,TESTED"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_INVA, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; -- skip header

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_A, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT("FAILURE! invalid assignment to INPUT_A");

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_ENA);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_B);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_ENB);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_F);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_CARRY_IN);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_CARRY_OUT);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_OUTPUT);

            INVA <= INPUT_INVA;
            A <= INPUT_A;
            ENA <= INPUT_ENA;
            B <= INPUT_B;
            ENB <= INPUT_ENB;
            F <= INPUT_F;
            CARRY_IN <= INPUT_CARRY_IN;
            CARRY_OUT_EXPECT <= INPUT_CARRY_OUT;
            OUTPUT_EXPECT <= INPUT_OUTPUT;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, INVA);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, A);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, ENA);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, B);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, ENB);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, F);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_IN);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_OUT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_OUT_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, OUTPUT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, OUTPUT_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            IF (CARRY_OUT = CARRY_OUT_EXPECT AND OUTPUT = OUTPUT_EXPECT) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;

        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;

    END PROCESS;
END TB;
