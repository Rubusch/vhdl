LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- port : the pinout for the modul
ENTITY BLINKY_ENT IS
PORT( BLINKY_CLK_50 : IN STD_LOGIC
 	; BLINKY_LED    : OUT STD_LOGIC := '0'
);
END ENTITY BLINKY_ENT;

-- architecture: the behavior implementation
ARCHITECTURE BLINKY_ARCH OF BLINKY_ENT IS
	SIGNAL HPS_RESET_N : STD_LOGIC;

	-- MACRO USING PRAGMA TRICK: FOR SETTING DIFFERENT VALUES FOR SIM AND SYNTH
	FUNCTION CLOCK_FREQUENCY RETURN NATURAL IS
	BEGIN
		-- SYNTHESIS TRANSLATE_OFF
		RETURN 50;
		-- SYNTHESIS TRANSLATE_ON
		RETURN 50000000;
	END CLOCK_FREQUENCY;

	CONSTANT CLK_FRQ : INTEGER := CLOCK_FREQUENCY;

BEGIN

	P1 : PROCESS(BLINKY_CLK_50, HPS_RESET_N)
		VARIABLE COUNTER : INTEGER := 0;
	BEGIN
        -- on top level check for event in respect to the above sensivity list
		IF HPS_RESET_N = '1' THEN
            -- try to always handle async reset events in a serializable manner
			COUNTER := 0;
		ELSIF RISING_EDGE(BLINKY_CLK_50) THEN
            -- the actual behavior driven by clock edges
			COUNTER := COUNTER + 1;
			IF COUNTER < CLK_FRQ THEN
				BLINKY_LED <= '1';
			ELSIF COUNTER >= CLK_FRQ AND COUNTER < 2*CLK_FRQ THEN
				BLINKY_LED <= '0';
			ELSE
				COUNTER := 0;
			END IF;
		END IF;
	END PROCESS P1;

END ARCHITECTURE BLINKY_ARCH;
