-- de1soc: adaptation for hardware
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_MODCOUNTER IS
GENERIC( MODULO : INTEGER := 16
    ; NBITS : INTEGER := 4
);
PORT( CLK50 : IN STD_LOGIC
    ; KEY_RST : IN STD_LOGIC
    ; HEX0_SEG : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    ; LED_COMPLETE_TICK : OUT STD_LOGIC
);
END DE1SOC_MODCOUNTER;

ARCHITECTURE DE1SOC OF DE1SOC_MODCOUNTER IS
    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';
    SIGNAL COMPLETE_TICK : STD_LOGIC := '0';
    SIGNAL COUNT : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0) := (OTHERS => '0');

    SIGNAL DATA : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL SEG : STD_LOGIC_VECTOR(6 DOWNTO 0) := (OTHERS => '0');

    SIGNAL PULSE : STD_LOGIC := '0';
    SIGNAL CLK_SCALED : STD_LOGIC := '0';

BEGIN

    FSMODCOUNTER : ENTITY WORK.FSMODCOUNTER
        GENERIC MAP (NBITS => NBITS, MODULO => MODULO)
        PORT MAP (CLK => CLK_SCALED, RST => RST, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

    SEVENSEG_UNIT : ENTITY WORK.DE1SOC_SEVENSEG
        PORT MAP (DATA => DATA, SEG => SEG);

    CLOCKSCALER_UNIT : ENTITY WORK.CLOCKSCALER
        GENERIC MAP (MODULO => 50000000, NBITS => 26)
        PORT MAP (CLK => CLK, RST => RST, PULSE => PULSE);

    -- WIRERING: IN
    CLK <= CLK50;
    RST <= NOT KEY_RST;

    -- WIRERING
    DATA <= COUNT;
    CLK_SCALED <= PULSE;

    -- WIRERIGN: OUT
    HEX0_SEG <= SEG;
    LED_COMPLETE_TICK <= COMPLETE_TICK;

END DE1SOC;
