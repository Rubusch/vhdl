-- hw adaptation for DE1SoC Board: dregister
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_DREGISTER IS
GENERIC( NBITS : INTEGER := 8 );
PORT( CLK50 : IN STD_LOGIC
    ; KEY : IN STD_LOGIC
    ; SW_ENA : IN STD_LOGIC)
    ; SW : IN STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
    ; LED : OUT STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
END DE1SOC_DREGISTER;

ARCHITECTURE DE1SOC OF DE1SOC_DREGISTER IS
    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';
    SIGNAL ENA : STD_LOGIC := '0';
    SIGNAL D : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL Q : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0) := (OTHERS => '0');

BEGIN

    DREGISTER_UNIT : ENTITY WORK.DREGISTER
        PORT MAP (CLK => CLK, RST => RST, ENA => ENA, D => D, Q => Q);

    -- IN
    CLK <= CLK50;
    RST <= NOT KEY;
    ENA <= SW_ENA;
    D <= SW;

    -- OUT
    LED <= Q;
END DE1SOC;
