-- hw adapter: full-adder
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_FULLADDER IS
PORT( SW_A : IN STD_LOGIC
    ; SW_B : IN STD_LOGIC
    ; SW_CARRY_IN : IN STD_LOGIC
    ; LED_SUM : OUT STD_LOGIC
    ; LED_CARRY_OUT : OUT STD_LOGIC
);
END DE1SOC_FULLADDER;

ARCHITECTURE DE1SOC OF DE1SOC_FULLADDER IS
    SIGNAL A : STD_LOGIC := '0';
    SIGNAL B : STD_LOGIC := '0';
    SIGNAL CARRY_IN : STD_LOGIC := '0';
    SIGNAL SUM : STD_LOGIC := '0';
    SIGNAL CARRY_OUT : STD_LOGIC := '0';

BEGIN

    FULLADDER_UNIT : ENTITY WORK.FULLADDER
        PORT MAP (A => A, B => B, CARRY_IN => CARRY_IN, SUM => SUM, CARRY_OUT => CARRY_OUT);

    -- IN
    A <= SW_A;
    B <= SW_B;
    CARRY_IN <= SW_CARRY_IN;

    -- OUT
    LED_SUM <= SUM;
    LED_CARRY_OUT <= CARRY_OUT;
END DE1SOC;
