--
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY MODCOUNTER_TB IS
END MODCOUNTER_TB;

ARCHITECTURE TB OF MODCOUNTER_TB IS
    CONSTANT T : TIME := 20 NS;
    -- TODO
BEGIN
    -- TODO
END TB;
