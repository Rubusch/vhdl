-- de1soc: hw adaptation of lfsr
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DE1SOC_LFSR IS
GENERIC( NBITS : INTEGER := 3);
PORT( CLK50 : IN STD_LOGIC
    ; KEY_RST : IN STD_LOGIC
    ; LED_Q : OUT STD_LOGIC_VECTOR(NBITS DOWNTO 0)
);

ARCHITECTURE DE1SOC OF DE1SOC_LFSR IS
    SIGNAL PULSE : STD_LOGIC;
    SIGNAL CLK : STD_LOGIC;
    SIGNAL RST : STD_LOGIC;

BEGIN

    CLK <= PULSE;
    RST <= NOT KEY_RST;

    CLOCKSCALER_UNIT : ENTITY WORK.CLOCKSCALER
        GENERIC MAP (MODULO => 50000000, NBITS => 26)
        PORT MAP (CLK => CLK50, RST => RST, PULSE => PULSE);

    LFSR_UNIT : ENTITY WORK.LFSR
        GENERIC MAP (NBITS => NBITS)
        PORT MAP (CLK => CLK, RST = RST, Q => LED_Q);
END DE1SOC;
