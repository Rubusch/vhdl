--
-- FULL-ADDER FOR ALU
--

-- TODO