--
-- A SIMPLE D-FLIPFLOP DEMO
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFLIPFLOP_ENT IS
PORT( CLK : IN STD_LOGIC
	; D : IN STD_LOGIC
	; Q : OUT STD_LOGIC
	; QBAR : OUT STD_LOGIC
);
END ENTITY DFLIPFLOP_ENT;

ARCHITECTURE DFLIPFLOP_ARCH OF DFLIPFLOP_ENT IS

BEGIN

END ARCHITECTURE DFLIPFLOP_ARCH;
