--
--
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY COUNTER_TB IS
END COUNTER_TB;

ARCHITECTURE TB OF COUNTER_TB IS
    CONSTANT T : TIME := 20 NS;
    SIGNAL CLK : STD_LOGIC;
    SIGNAL RST : STD_LOGIC;
    SIGNAL COMPLETE_TICK : STD_LOGIC;
    SIGNAL COUNT : STD_LOGIC_VECTOR(2 DOWNTO 0);

    CONSTANT NUM_OF_CLOCKS := 30;
    SIGNAL I : INTEGER := 0;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    COUNTER_UNIT : ENTITY WORK.COUNTER
        GENERIC MAP (N => '3')
        PORT MAP (CLK => CLK, RST => RST, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

-- TODO

END TB;
