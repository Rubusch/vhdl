--
-- LOGICAL UNIT FOR ALU
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LOGICAL_ENT IS
PORT( A : IN STD_LOGIC
    ; B : IN STD_LOGIC
    ; SELECT_AND : IN STD_LOGIC
    ; SELECT_OR : IN STD_LOGIC
    ; SELECT_NOT : IN STD_LOGIC
    ; OUTPUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END ENTITY LOGICAL_ENT;

ARCHITECTURE LOGICAL_ARCH OF LOGICAL_ENT IS
    SIGNAL A_AND_B : STD_LOGIC;
    SIGNAL A_OR_B : STD_LOGIC;
    SIGNAL NOT_B : STD_LOGIC;
BEGIN
    A_AND_B <= SELECT_AND AND (A AND B);
    A_OR_B <= SELECT_OR AND (A OR B);
    NOT_B <= SELECT_NOT AND (NOT B);

    OUTPUT <= (A_AND_B, A_OR_B, NOT_B);
--    OUTPUT <= STD_LOGIC_VECTOR(NOT_B, A_OR_B, A_AND_B); -- TODO TEST WHICH ONE TO TAKE?
END ARCHITECTURE LOGICAL_ARCH;
