-- hw adaptation for DE1SoC board (cycloneV)
--
-- author: Lothar Rubusch

LIBARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_COUNTER IS
PORT( SW_D : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
    ; KEY_C : IN STD_LOGIC
    ; LED_S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END DE1SOC_COUNTER;

ARCHITECTURE DE1SOC OF DE1SOC_COUNTER IS
    SIGNAL D : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL C : STD_LOGIC;
    SIGNAL S : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

    COUNTER_UNIT : ENTITY WORK.COUNTER
        PORT MAP (D => D, C => C, S => S);

    -- IN
    D <= SW_D;
    C <= NOT KEY_C;

    -- OUT
    LED_S <= S;
END DE1SOC;
