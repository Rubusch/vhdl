-- tb: decoder
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_DECODER IS
END TB_DECODER;

ARCHITECTURE TB OF TB_DECODER IS

BEGIN

END TB;
