-- tb: multiplexer
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_MULTIPLEXER IS
END TB_MULTIPLEXER;

ARCHITECTURE TB OF TB_MULTIPLEXER IS
    CONSTANT NBIT : INTEGER := 4;
    SIGNAL A : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL B : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL SEL : STD_LOGIC := '0';
    SIGNAL C : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL C_EXPECT : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    QUADMUX_UNIT : ENTITY WORK.QUADMUX
        GENERIC MAP (NBIT => NBIT)
        PORT MAP (A => A, B => B, SEL => SEL, C => C);

    PROCESS
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE GOOD_NUM : BOOLEAN;
        VARIABLE SEPARATOR : CHARACTER;
        VARIABLE INPUT_A : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
        VARIABLE INPUT_B : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
        VARIABLE INPUT_SEL : STD_LOGIC;
        VARIABLE INPUT_C : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("A,B,SEL,C,C_EXPECT,TESTED"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_A, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM;

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_B, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT("FAILURE! invalid assignment to INPUT_B");

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_SEL);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_C);

            A <= INPUT_A;
            B <= INPUT_B;
            SEL <= INPUT_SEL;
            C_EXPECT <= INPUT_C;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, A);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, B);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, SEL);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, C);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, C_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            IF (C = C_EXPECT) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;
        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;
    END PROCESS;
END TB;
