-- mod counter as state machine
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FSMCOUNTER IS
GENERIC( MODULO : NATURAL := 6
    ; NBITS : NATURAL := 4
);
PORT( CLK : IN STD_LOGIC
    ; RST : IN STD_LOGIC
    ; OUT_MOORE : OUT STD_LOGIC_VECTOR(NBITES-1 DOWNTO 0);
);
END FSMCOUNTER;

ARCHITECTURE FSM OF FSMCOUNTER IS
    TYPE STATETYPE_MOORE (START_MOORE, COUNT_MOORE);
    SIGNAL STATE_MOORE_REG, STATE_MOORE_NEXT : STATETYPE_MOORE;
    SIGNAL COUNT_MOORE_REG, COUNT_MOORE_NEXT : UNSIGNED(NBITS-1 DOWNTO 0);

BEGIN

    PROCESS(CLK, RST)
    BEGIN
        IF (RST = '1') THEN
            STATE_MOORE_REG <= START_MOORE;
            COUNT_MOORE_REG <= (OTHERS => '0');
        ELSIF (RISING_EDGE(CLK)) THEN
            STATE_MOORE_REG <= STATE_MOORE_NEXT;
            COUNT_MOORE_REG <= COUNT_MOORE_NEXT;
        END IF;
    END PROCESS;

    PROCESS(COUNT_MOORE_REG, STATE_MOORE_REG)
    BEGIN
        CASE STATE_MOORE_REG IS
            WHEN START_MOORE =>
                COUNT_MOORE_NEXT <= (OTHERS => '0');
                STATE_MOORE_NEXT <= COUNT_MOORE;
            WHEN COUNT_MODE =>
                COUNT_MOORE_NEXT <= COUNT_MOORE_REG + 1;
                IF ((COUNT_MOORE_REG + 1) = MODULO -1) THEN
                    STATE_MOORE_NEXT <= START_MOORE;
                ELSE
                    STATE_MOORE_NEXT <= COUNT_MOORE;
                END IF;
        END CASE;
    END PROCESS;

    OUT_MOORE <= STD_LOGIC_VECTOR(COUNT_MOORE_REG);
END FSM
