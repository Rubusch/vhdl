-- tb: glitch02
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_GLITCHY IS
END TB_GLITCHY;

ARCHITECTURE TB OF TB_GLITCHY IS
    CONSTANT T : TIME := 20 NS;
    CONSTANT NCLKS : INTEGER := 50;
    SIGNAL I : INTEGER := 0;

    FILE OUTPUT_BUF : TEXT;

    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL DIN : STD_LOGIC := '0';
    SIGNAL DOUT : STD_LOGIC := '0';

BEGIN

    GLITCHY_UNIT : ENTITY WORK.GLITCHY
        PORT MAP (CLK => CLK, DIN => DIN, DOUT => DOUT);

    PROCESS
    BEGIN
        CLK <= '0';
        WAIT FOR T/2;
        CLK <= '1';
        WAIT FOR T/2;
        IF (I = NCLKS) THEN
            FILE_CLOSE(OUTPUT_BUF);
            WAIT;
        ELSE
            I <= I + 1;
        END IF;

        IF (I > 3 AND i < 6) THEN
            DIN <= '1';
        ELSE
            DIN <= '0';
        END IF;
    END PROCESS;

    FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

    PROCESS(CLK)
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
    BEGIN
        IF (CLK'EVENT AND CLK = '1') THEN
            IF (I = 0) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("CLK,DIN,DOUT"));
                WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
            END IF;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, CLK);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, DIN);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, DOUT);
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END IF;
    END PROCESS;
END TB;
