-- counter adaptation for DE1SoC Board
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_MODCOUNTER IS
GENERIC( NBITS : INTEGER := 2
    ; MAX_NUM : INTEGER := 4
);
PORT( CLK50 : IN STD_LOGIC
    ; KEY : IN STD_LOGIC
    ; LED : OUT STD_LOGIC
    ; LEDR : OUT STD_LOGIC_VECTOR()
);
END DE1SOC_MODCOUNTER;

ARCHITECTURE HW OF DE1SOC_MODCOUNTER IS
-- TODO
BEGIN
-- TODO
END HW;
