-- counter adaptation for DE1SoC Board
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_MODCOUNTER IS
-- TODO
END DE1SOC_MODCOUNTER;

ARCHITECTURE HW OF DE1SOC_MODCOUNTER IS
-- TODO
BEGIN
-- TODO
END HW;
