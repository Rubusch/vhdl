LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DREGISTER_ENT IS
PORT( D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    CLK : IN STD_LOGIC;
    ENA : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    Q   : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
END ENTITY DREGISTER_ENT;


