--
-- FULL-ADDER FOR ALU
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FULLADDER IS
PORT( A : IN STD_LOGIC
    ; B : IN STD_LOGIC
    ; CARRY_IN : IN STD_LOGIC
    ; CARRY_OUT : OUT STD_LOGIC
    ; SUM : OUT STD_LOGIC
    ; SEL : IN STD_LOGIC
);
END ENTITY FULLADDER;

ARCHITECTURE FULLADDER_ARCH OF FULLADDER IS
    SIGNAL SUM_TMP : STD_LOGIC := '0';
BEGIN
    SUM_TMP <= A XOR B;
    CARRY_OUT <= (SEL AND A AND B) OR (SEL AND SUM_TMP AND CARRY_IN);
    SUM <= SEL AND (CARRY_IN XOR SUM_TMP);
END ARCHITECTURE FULLADDER_ARCH;
