--
-- DECODER FOR ALU
--

-- TODO