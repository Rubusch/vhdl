--
-- LOGICAL UNIT FOR ALU
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LOGICAL_ENT IS
PORT( A : IN STD_LOGIC
    ; B : IN STD_LOGIC
    ; SELECT_AND : IN STD_LOGIC
    ; SELECT_OR : IN STD_LOGIC
    ; SELECT_NOT : IN STD_LOGIC
    ; OUTPUT : OUT STD_LOGIC
);
END ENTITY LOGICAL_ENT;

ARCHITECTURE LOGICAL_ARCH OF LOGICAL_ENT IS
    SIGNAL A_AND_B : STD_LOGIC;
    SIGNAL A_OR_B : STD_LOGIC;
    SIGNAL NOT_B : STD_LOGIC;
BEGIN
    A_AND_B <= SELECT_AND AND (A AND B);
    A_OR_B <= SELECT_OR AND (A OR B);
    NOT_B <= SELECT_NOT AND (NOT B);

    OUTPUT <= A_AND_B OR A_OR_B OR NOT_B;
END ARCHITECTURE LOGICAL_ARCH;
