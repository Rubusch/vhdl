-- mod counter as state machine
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FSMCOUNTER IS
GENERIC( MODULO : NATURAL := 6
    ; NBITS : NATURAL := 4
);
PORT( CLK : IN STD_LOGIC
    ; RST : IN STD_LOGIC
    ; COMPLETE_TICK : OUT STD_LOGIC
    ; COUNT : OUT STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
);
END FSMCOUNTER;

ARCHITECTURE FSM OF FSMCOUNTER IS
    SIGNAL COUNT_MOORE_REG, COUNT_MOORE_NEXT : UNSIGNED(NBITS-1 DOWNTO 0);
    TYPE STATETYPE_MOORE IS (START_MOORE, COUNT_MOORE);
    SIGNAL STATE_MOORE_REG, STATE_MOORE_NEXT : STATETYPE_MOORE;

BEGIN

    PROCESS(CLK, RST)
    BEGIN
        IF (RST = '1') THEN
            COUNT_MOORE_REG <= (OTHERS => '0');
            STATE_MOORE_REG <= START_MOORE;
        ELSIF (RISING_EDGE(CLK)) THEN
            COUNT_MOORE_REG <= COUNT_MOORE_NEXT;
            STATE_MOORE_REG <= STATE_MOORE_NEXT;
        END IF;
        COUNT <= STD_LOGIC_VECTOR(COUNT_MOORE_REG);
    END PROCESS;

    PROCESS(COUNT_MOORE_REG, STATE_MOORE_REG)
    BEGIN
        CASE STATE_MOORE_REG IS
            WHEN START_MOORE =>
                COUNT_MOORE_NEXT <= (OTHERS => '0');
                STATE_MOORE_NEXT <= COUNT_MOORE;
                COMPLETE_TICK <= '0';
            WHEN COUNT_MOORE =>
                COUNT_MOORE_NEXT <= COUNT_MOORE_REG + 1;
                IF ((COUNT_MOORE_REG + 1) = MODULO - 1) THEN
                    COMPLETE_TICK <= '1';
                    STATE_MOORE_NEXT <= START_MOORE;
                ELSE
                    COMPLETE_TICK <= '0';
                    STATE_MOORE_NEXT <= COUNT_MOORE;
                END IF;
        END CASE;
    END PROCESS;

END FSM;
