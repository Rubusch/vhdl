-- hw adaptation: comparator
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_COMPARATOR IS
PORT( SW_A : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; SW_B : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; LED_Q : OUT STD_LOGIC
);
END DE1SOC_COMPARATOR;

ARCHITECTURE DE1SOC OF DE1SOC_COMPARATOR IS
    SIGNAL A : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL B : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL Q : STD_LOGIC := '0';

BEGIN

    COMPARATOR_UNIT : ENTITY WORK.COMPARATOR
        PORT MAP (A => A, B => B, Q => Q);

    -- IN
    A <= SW_A;
    B <= SW_B;

    -- OUT
    LED_Q <= Q;
END DE1SOC;
