-- testbench: andnand
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_ANDNAND IS
END TB_ANDNAND;

ARCHITECTURE TB OF TB_ANDNAND IS
    SIGNAL A : STD_LOGIC;
    SIGNAL B : STD_LOGIC;
    SIGNAL Q : STD_LOGIC;
    SIGNAL Q_EXPECT : STD_LOGIC;
    SIGNAL QBAR : STD_LOGIC;
    SIGNAL QBAR_EXPECT : STD_LOGIC;

    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    ANDNAND_UNIT : ENTITY WORK.ANDNAND
        PORT MAP (A => A, B => B, Q => Q, QBAR => QBAR);

    PROCESS
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE INPUT_A : STD_LOGIC;
        VARIABLE INPUT_B : STD_LOGIC;
        VARIABLE INPUT_Q : STD_LOGIC;
        VARIABLE INPUT_QBAR : STD_LOGIC;
        VARIABLE SEPARATOR : CHARACTER;
        VARIABLE GOOD_NUM ; BOOLEAN;
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("A,B,Q,Q_EXPECT,QBAR,QBAR_EXPECT"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            -- header
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_A, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; -- skip head line

            -- read input
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_B, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT "FAILURE! bad value for B";

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_Q);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_QBAR);

            A <= INPUT_A;
            B <= INPUT_B;
            Q_EXPECT <= INPUT_Q;
            QBAR_EXPECT <= INPUT_QBAR;

            -- execute
            WAIT FOR 20 NS;

            -- write results
            WRITE(WRITE_COL_TO_OUTPUT_BUF, A);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, B);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, Q);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, Q_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, QBAR);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, QBAR_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            IF ((Q = Q_EXPECT) AND (QBAR = QBAR_EXPECT)) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;

        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;

    END PROCESS;
END TB;

