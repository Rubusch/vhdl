--
--
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY COUNTER_TB IS
END COUNTER_TB;

ARCHITECTURE TB OF COUNTER_TB IS
    CONSTANT T : TIME := 20 NS;
    SIGNAL CLK : STD_LOGIC;
    SIGNAL RST : STD_LOGIC;
    SIGNAL COMPLETE_TICK : STD_LOGIC;
    SIGNAL COUNT : STD_LOGIC_VECTOR(2 DOWNTO 0);

    CONSTANT NUM_OF_CLOCKS : INTEGER := 30; -- TODO test
    SIGNAL I : INTEGER := 0;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    COUNTER_UNIT : ENTITY WORK.COUNTER
        GENERIC MAP (N => '3')
        PORT MAP (CLK => CLK, RST => RST, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

    RST <= '1', '0' AFTER T/2;

    PROCESS
    BEGIN
        CLK <= '0';
        WAIT FOR T/2;
        CLK <= '1';
        WAIT FOR T/2;
        IF (I = NUM_OF_CLOCKS) THEN
            FILE_CLOSE(OUTPUT_BUF);
            WAIT;
        ELSE
            I <= I + 1;
        END IF;
    END PROCESS;

    FILE_OPEN(OUTPUT_BUF, "../../results_tb.csv", WRITE_MODE);

    PROCESS(CLK)
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
    BEGIN
        IF (CLK'EVENT AND CLK = '1' AND RST /= '1') THEN
            IF (I = '0') THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("RST,COMPLETE_TICK,COUNT"));
                WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
            END IF;
            WRITE(WRITE_COL_TO_OUTPUT_BUF, RST);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, COMPLETE_TICK);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, COUNT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END IF;
    END PROCESS;
END TB;
