-- MODMCOUNTER_TB.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MODMCOUNTER_ENT_TB IS
END MODMCOUNTER_ENT_TB;

ARCHITECTURE TB OF MODMCOUNTER_ENT_TB IS
    CONSTANT M : INTEGER := 10;
    CONSTANT N : INTEGER := 4;
    CONSTANT T : TIME := 20 NS;

    SIGNAL CLK, RESET : STD_LOGIC; -- input
    SIGNAL COMPLETE_TICK : STD_LOGIC; -- output
    SIGNAL COUNT : STD_LOGIC_VECTOR(N-1 DOWNTO 0); -- output

BEGIN

    MODMCOUNTER_UNIT : ENTITY WORK.MODMCOUNTER_ENT
        GENERIC MAP (M => M, N => N)
        PORT MAP (CLK => CLK, RESET => RESET, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

    -- continuous clock
    PROCESS
    BEGIN
        CLK <= '0';
        WAIT FOR T/2;
        CLK <= '1';
        WAIT FOR T/2;
    END PROCESS;

    -- reset = 1 for first clock cycle, then 0
    RESET <= '1', '0' AFTER T/2;
END TB;
