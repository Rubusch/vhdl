-- hw adaptation for DE1SoC Board: d-flipflop
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_DFLIPFLOP IS
PORT( CLK50, KEY, SW : IN STD_LOGIC
    ; LED : OUT STD_LOGIC
);
END DE1SOC_DFLIPFLOP;

ARCHITECTURE HW OF DE1SOC_DFLIPFLOP IS
    SIGNAL CLK, RST, D, Q : STD_LOGIC;

BEGIN

    DFLIPFLOP_UNIT : ENTITY WORK.DFLIPFLOP
        PORT MAP (CLK => CLK, RST => RST, D => D, Q => Q);

    -- IN
    CLK <= CLK50;
    RST <= NOT KEY;
    D <= SW;

    -- OUT
    LED <= Q;
END HW;
