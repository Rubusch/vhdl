-- tb: mealy and moore
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_MEALYANDMOORE IS
END TB_MEALYANDMOORE;

ARCHITECTURE TB OF TB_MEALYANDMOORE IS
    CONSTANT T : TIME := 20 NS;
    CONSTANT NCLKS : INTEGER := 50;
    SIGNAL I : INTEGER := 0;

    FILE OUTPUT_BUF : TEXT;

    SIGNAL MEALY_TICK : STD_LOGIC := '0';
    SIGNAL MOORE_TICK : STD_LOGIC := '0';
    SIGNAL LEVEL : STD_LOGIC := '0';

    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';

BEGIN

    MEALYANDMOORE_UNIT : ENTITY WORK.MEALYANDMOORE
        PORT MAP (CLK => CLK, RST => RST, LEVEL => LEVEL, MEALY_TICK => MEALY_TICK, MOORE_TICK => MOORE_TICK);

    RST <= '1', '0' AFTER T/2;

    PROCESS
    BEGIN
        CLK <= '0';
        WAIT FOR T/2;
        CLK <= '1';
        WAIT FOR T/2;
        IF (I = NCLKS) THEN
            FILE_CLOSE(OUTPUT_BUF);
            WAIT;
        ELSE
            I <= I + 1;
        END IF;

        IF (I > 2 AND I < 6) THEN
            LEVEL <= '1';
        ELSE
            LEVEL <= '0';
        END IF;
    END PROCESS;

    FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

    PROCESS(CLK)
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
    BEGIN
        IF (CLK'EVENT AND CLK = '1' AND RST /= '1') THEN
            IF (I = 0) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("LEVEL,MEALY_TICK,MOORE_TICK"));
                WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
            END IF;
            WRITE(WRITE_COL_TO_OUTPUT_BUF, LEVEL);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, MEALY_TICK);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, MOORE_TICK);
            
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END IF;
    END PROCESS;
END TB;
