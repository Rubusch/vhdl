-- testscreen: display four squares of different color on the screen
--
-- author: Lothar Rubusch
-- original from: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_TESTSCREEN IS
GENERIC( PIXEL_WIDTH : INTEGER := 10 );
PORT( CLK : IN STD_LOGIC
    ; RST : IN STD_LOGIC
    ; VGA_CLK : OUT STD_LOGIC
    ; VGA_BLANK_N : OUT STD_LOGIC
    ; VGA_HS : OUT STD_LOGIC
    ; VGA_VS : OUT STD_LOGIC
    ; VGA_R : OUT STD_LOGIC_VECTOR(PIXEL_WIDTH-1 DOWNTO 0)
    ; VGA_G : OUT STD_LOGIC_VECTOR(PIXEL_WIDTH-1 DOWNTO 0)
    ; VGA_B : OUT STD_LOGIC_VECTOR(PIXEL_WIDTH-1 DOWNTO 0)
);
END DE1SOC_TESTSCREEN;

ARCHITECTURE DE1SOC OF DE1SOC_TESTSCREEN IS
    SIGNAL RGB_REG : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
    SIGNAL VIDEO_ON : STD_LOGIC := '0';
    SIGNAL PIXEL_X : STD_LOGIC_VECTOR(PIXEL_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL PIXEL_Y : STD_LOGIC_VECTOR(PIXEL_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL PIX_X : INTEGER := 0;
    SIGNAL PIX_Y : INTEGER := 0;

BEGIN

END DE1SOC;
