LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BLINKY_ENT IS
PORT    (BLINKY_CLK_50 : IN STD_LOGIC
 	;BLINKY_RST_N  : IN STD_LOGIC := '0'
 	;BLINKY_LED    : OUT STD_LOGIC
);
END ENTITY BLINKY_ENT;

ARCHITECTURE BLINKY_ARCH OF BLINKY_ENT IS
	-- MACRO USING PRAGMA TRICK: FOR SETTING DIFFERENT VALUES FOR SIM AND SYNTH
	FUNCTION CLOCK_FREQUENCY RETURN NATURAL IS
	BEGIN
		-- SYNTHESIS TRANSLATE_OFF
		RETURN 50;
		-- SYNTHESIS TRANSLATE_ON
		RETURN 50000000;
	END CLOCK_FREQUENCY;

	CONSTANT CLK_FRQ : INTEGER := CLOCK_FREQUENCY;

BEGIN

	P1 : PROCESS(BLINKY_CLK_50, BLINKY_RST_N)
	VARIABLE COUNTER : INTEGER := 0;
	BEGIN
		IF BLINKY_RST_N = '1' THEN
			COUNTER := 0;
		ELSIF RISING_EDGE(BLINKY_CLK_50) THEN
			COUNTER := COUNTER + 1;
			IF COUNTER < CLK_FRQ THEN
				BLINKY_LED <= '1';
			ELSIF COUNTER >= CLK_FRQ THEN
				BLINKY_LED <= '0';
			ELSE
--			BLINKY_LED <= (COUNTER < CLK_FRQ);
--			IF COUNTER > 2*CLK_FRQ THEN
				COUNTER := 0;
			END IF;
		END IF;
	END PROCESS P1;

END ARCHITECTURE BLINKY_ARCH;
