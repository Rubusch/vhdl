-- half-adder_tb.vhd

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY FULLADDER_TB IS
END FULLADDER_TB;

ARCHITECTURE TB OF FULLADDER_TB IS
    SIGNAL A, B, CARRY_IN : STD_LOGIC;
    SIGNAL SUM_EXPECTED, CARRY_OUT_EXPECTED : STD_LOGIC;
    SIGNAL SUM, CARRY_OUT : STD_LOGIC;
    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    CONNECTION : ENTITY WORK.fulladder PORT MAP (
        A => A,
        B => B,
        CARRY_IN => CARRY_IN,
        SUM => SUM,
        CARRY_OUT => CARRY_OUT);

    TB1 : PROCESS
    VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
    VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
    VARIABLE VAL_A, VAL_B, VAL_CARRY_IN : STD_LOGIC;
    VARIABLE VAL_SUM, VAL_CARRY_OUT : STD_LOGIC;
    VARIABLE VAL_SEPARATOR : CHARACTER;
    VARIABLE GOOD_NUM : BOOLEAN;
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../result.csv", WRITE_MODE);
        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("A,B,CARRY_IN,SUM,SUM_EXPECTED,CARRY_OUT,CARRY_OUT_EXPECTED,RESULT"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, VAL_A, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; -- i.e. skip the header line

            READ(READ_COL_FROM_INPUT_BUF, VAL_SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, VAL_B, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT "BAD VALUE ASSIGNED TO VAL_B";

            READ(READ_COL_FROM_INPUT_BUF, VAL_SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, VAL_CARRY_IN);
            READ(READ_COL_FROM_INPUT_BUF, VAL_SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, VAL_SUM);
            READ(READ_COL_FROM_INPUT_BUF, VAL_SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, VAL_CARRY_OUT);

            A <= VAL_A;
            B <= VAL_B;
            CARRY_IN <= VAL_CARRY_IN;
            SUM_EXPECTED <= VAL_SUM;
            CARRY_OUT_EXPECTED <= VAL_CARRY_OUT;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, A);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, B);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_IN);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, SUM);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, SUM_EXPECTED);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_OUT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, CARRY_OUT_EXPECTED);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));

            IF ((SUM_EXPECTED = SUM) AND (CARRY_OUT_EXPECTED = CARRY_OUT)) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK,"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL,"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;

        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;

    END PROCESS;
END TB;
