--
-- FULL-ADDER FOR ALU
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FULLADDER_ENT IS
PORT( A : IN STD_LOGIC
    ; B : IN STD_LOGIC
    ; CARRY_IN : IN STD_LOGIC
    ; CARRY_OUT : OUT STD_LOGIC
    ; SUM : OUT STD_LOGIC
    ; SEL : IN STD_LOGIC
);
END ENTITY FULLADDER_ENT;

ARCHITECTURE FULLADDER_ARCH OF FULLADDER_ENT IS
    SIGNAL SUM_TMP : STD_LOGIC;
BEGIN
    SUM_TMP <= A XOR B;
    CARRY_OUT <= (SEL AND A AND B) OR (SEL AND SUM_TMP AND CARRY_IN);
    SUM <= SEL AND (CARRY_IN XOR SUM_TMP);
END ARCHITECTURE FULLADDER_ARCH;
