-- tb: clockscaler
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_CLOCKSCALER IS
END TB_CLOCKSCALER;

ARCHITECTURE TB OF TB_CLOCKSCALER IS
    

BEGIN

    CLOCKSCALER_UNIT : ENTITY WORK.CLOCKSCALER 
        PORT MAP
END TB;
