--
--
--
--
--
--
--
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DECORATOR_ENT IS
PORT( A : IN STD_LOGIC := '0'
    ; B : IN STD_LOGIC := '0'
    ; C : IN STD_LOGIC := '0'
    ; D : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ENTITY DECORATOR_ENT;

ARCHITECTURE DECORATOR_ARCH OF DECORATOR_ENT IS

BEGIN

END ARCHITECTURE DECORATOR_ARCH;
