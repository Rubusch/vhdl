-- tb: shifter
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_SHIFTER IS
END TB_SHIFTER;

ARCHITECTURE TB OF TB_SHIFTER IS
    SIGNAL D : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    SIGNAL C : STD_LOGIC := '0';
    SIGNAL S : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    SIGNAL S_EXPECT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    SHIFTER_UNIT : ENTITY WORK.SHIFTER
        PORT MAP (D => D, C => C, S => S);

    PROCESS
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE GOOD_NUM : BOOLEAN;
        VARIABLE SEPARATOR : CHARACTER;
        VARIABLE INPUT_D : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
        VARIABLE INPUT_C : STD_LOGIC := '0';
        VARIABLE INPUT_S : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("D,C,S,S_EXPECT,TESTED"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_D, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; -- skip header

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_C, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT "FAILURE! bad value assigned to D";

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_S);

            D <= INPUT_D;
            C <= INPUT_C;
            S_EXPECT <= INPUT_S;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, D);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, C);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, S);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, S_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));

            IF (S = S_EXPECT) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;

        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;
    END PROCESS;
END TB;
