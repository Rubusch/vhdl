-- hw adaptation for DE1SoC Board: fsm
-- (visual verification)
--
-- Author: Lothar Rubusch

-- TODO
