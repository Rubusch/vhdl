--
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY MODCOUNTER_TB IS
END MODCOUNTER_TB;

ARCHITECTURE TB OF MODCOUNTER_TB IS
    CONSTANT T : TIME := 20 NS;
    CONSTANT NBITS : UNSIGNED := 2;
    CONSTANT MAX_NUM : UNSIGNED := 4;
    SIGNAL CLK : STD_LOGIC;
    SIGNAL RST : STD_LOGIC;
    SIGNAL COMPLETE_TICK : STD_LOGIC;
    SIGNAL COUNT : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0);

    CONSTANT NUM_OF_CLOCKS : INTEGER := 30;
    SIGNAL I : INTEGER := 0;

    FILE OUTPUT_BUF : TEXT;

BEGIN

    
    -- TODO
END TB;
