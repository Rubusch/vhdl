-- de1soc: hw adaptation for serial parallel converter via shifter
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

-- TODO
