-- de1soc: hw adapter for dual port ram
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_DUALPORTRAM IS
GENERIC( ADDR_WIDTH : INTEGER := 2
    ; DATA_WIDTH : INTEGER := 3
);
PORT( CLK50 : IN STD_LOGIC
    ; SW_WE : IN STD_LOGIC
    ; SW_ADDR_WR : IN STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0)
    ; SW_ADDR_RD : IN STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0)
    ; SW_DIN : IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
    ; LED_DOUT : OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
);
END DE1SOC_DUALPORTRAM;

ARCHITECTURE DE1SOC OF DE1SOC_DUALPORTRAM IS
BEGIN

    DUALPORTRAM_UNIT : ENTITY WORK.DUALPORTRAM
        PORT MAP (CLK => CLK50, WE => SW_WE, ADDR_WR => SW_ADDR_WR, ADDR_RD => SW_ADDR_RD, DIN => SW_DIN, DOUT => LED_DOUT);
END DE1SOC;
