// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Build 646 04/11/2019 SJ Lite Edition"

// DATE "08/24/2020 18:59:31"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module sdram_demo (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	led_export,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	sw_export)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
output 	[7:0] led_export;
output 	[12:0] sdram_wire_addr;
output 	[1:0] sdram_wire_ba;
output 	sdram_wire_cas_n;
output 	sdram_wire_cke;
output 	sdram_wire_cs_n;
inout 	[31:0] sdram_wire_dq;
output 	[3:0] sdram_wire_dqm;
output 	sdram_wire_ras_n;
output 	sdram_wire_we_n;
input 	[7:0] sw_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdram|m_addr[0]~q ;
wire \sdram|m_addr[1]~q ;
wire \sdram|m_addr[2]~q ;
wire \sdram|m_addr[3]~q ;
wire \sdram|m_addr[6]~q ;
wire \sdram|m_addr[7]~q ;
wire \sdram|m_addr[8]~q ;
wire \sdram|m_addr[9]~q ;
wire \nios2|cpu|W_alu_result[4]~q ;
wire \nios2|cpu|W_alu_result[5]~q ;
wire \nios2|cpu|W_alu_result[9]~q ;
wire \nios2|cpu|W_alu_result[24]~q ;
wire \nios2|cpu|W_alu_result[25]~q ;
wire \nios2|cpu|W_alu_result[26]~q ;
wire \nios2|cpu|W_alu_result[27]~q ;
wire \nios2|cpu|W_alu_result[28]~q ;
wire \nios2|cpu|W_alu_result[20]~q ;
wire \nios2|cpu|W_alu_result[19]~q ;
wire \nios2|cpu|W_alu_result[21]~q ;
wire \nios2|cpu|W_alu_result[22]~q ;
wire \nios2|cpu|W_alu_result[23]~q ;
wire \nios2|cpu|W_alu_result[18]~q ;
wire \nios2|cpu|W_alu_result[17]~q ;
wire \nios2|cpu|W_alu_result[16]~q ;
wire \nios2|cpu|W_alu_result[15]~q ;
wire \nios2|cpu|W_alu_result[14]~q ;
wire \nios2|cpu|W_alu_result[13]~q ;
wire \nios2|cpu|W_alu_result[6]~q ;
wire \nios2|cpu|W_alu_result[7]~q ;
wire \nios2|cpu|W_alu_result[8]~q ;
wire \nios2|cpu|W_alu_result[12]~q ;
wire \nios2|cpu|W_alu_result[11]~q ;
wire \nios2|cpu|W_alu_result[10]~q ;
wire \nios2|cpu|W_alu_result[2]~q ;
wire \nios2|cpu|W_alu_result[3]~q ;
wire \nios2|cpu|F_pc[17]~q ;
wire \nios2|cpu|F_pc[16]~q ;
wire \nios2|cpu|F_pc[18]~q ;
wire \nios2|cpu|F_pc[19]~q ;
wire \nios2|cpu|F_pc[20]~q ;
wire \nios2|cpu|F_pc[21]~q ;
wire \nios2|cpu|F_pc[22]~q ;
wire \nios2|cpu|F_pc[23]~q ;
wire \nios2|cpu|F_pc[24]~q ;
wire \nios2|cpu|F_pc[26]~q ;
wire \nios2|cpu|F_pc[15]~q ;
wire \nios2|cpu|F_pc[14]~q ;
wire \nios2|cpu|F_pc[9]~q ;
wire \nios2|cpu|F_pc[11]~q ;
wire \nios2|cpu|F_pc[13]~q ;
wire \nios2|cpu|F_pc[12]~q ;
wire \nios2|cpu|F_pc[10]~q ;
wire \nios2|cpu|F_pc[0]~q ;
wire \nios2|cpu|F_pc[1]~q ;
wire \nios2|cpu|F_pc[2]~q ;
wire \nios2|cpu|F_pc[3]~q ;
wire \nios2|cpu|F_pc[4]~q ;
wire \nios2|cpu|F_pc[5]~q ;
wire \nios2|cpu|F_pc[6]~q ;
wire \nios2|cpu|F_pc[7]~q ;
wire \nios2|cpu|F_pc[8]~q ;
wire \sdram|oe~q ;
wire \ram|the_altsyncram|auto_generated|ram_block1a32~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a0~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a54~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a22~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a55~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a23~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a56~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a24~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a57~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a25~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a58~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a26~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a33~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a1~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a36~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a4~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a35~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a3~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a34~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a2~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a43~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a11~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a44~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a12~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a45~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a13~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a46~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a14~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a47~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a15~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a48~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a16~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a37~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a5~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a40~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a8~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a42~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a10~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a41~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a9~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a60~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a28~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a53~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a21~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a61~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a29~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a62~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a30~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a63~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a31~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a49~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a17~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a50~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a18~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a59~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a27~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a39~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a7~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a38~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a6~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a52~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a20~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a51~portadataout ;
wire \ram|the_altsyncram|auto_generated|ram_block1a19~portadataout ;
wire \nios2|cpu|d_writedata[8]~q ;
wire \nios2|cpu|d_writedata[9]~q ;
wire \nios2|cpu|d_writedata[10]~q ;
wire \nios2|cpu|d_writedata[11]~q ;
wire \nios2|cpu|d_writedata[12]~q ;
wire \nios2|cpu|d_writedata[13]~q ;
wire \nios2|cpu|d_writedata[14]~q ;
wire \nios2|cpu|d_writedata[15]~q ;
wire \nios2|cpu|d_writedata[16]~q ;
wire \nios2|cpu|d_writedata[17]~q ;
wire \nios2|cpu|d_writedata[18]~q ;
wire \nios2|cpu|d_writedata[19]~q ;
wire \nios2|cpu|d_writedata[20]~q ;
wire \nios2|cpu|d_writedata[21]~q ;
wire \nios2|cpu|d_writedata[22]~q ;
wire \nios2|cpu|d_writedata[23]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[0]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[22]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[23]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[24]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[25]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[26]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[1]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[4]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[3]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[2]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[11]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[12]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[13]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[14]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[15]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[16]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[5]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[8]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[10]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[9]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[28]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[21]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[29]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[30]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[31]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[17]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[18]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[27]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[7]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[6]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[20]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[19]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \jtag_uart|Add1~1_sumout ;
wire \jtag_uart|Add1~5_sumout ;
wire \jtag_uart|Add1~9_sumout ;
wire \jtag_uart|Add1~13_sumout ;
wire \jtag_uart|Add1~17_sumout ;
wire \jtag_uart|Add1~21_sumout ;
wire \jtag_uart|Add1~25_sumout ;
wire \led|data_out[0]~q ;
wire \led|data_out[1]~q ;
wire \led|data_out[2]~q ;
wire \led|data_out[3]~q ;
wire \led|data_out[4]~q ;
wire \led|data_out[5]~q ;
wire \led|data_out[6]~q ;
wire \led|data_out[7]~q ;
wire \sdram|m_addr[4]~q ;
wire \sdram|m_addr[5]~q ;
wire \sdram|m_addr[10]~q ;
wire \sdram|m_addr[11]~q ;
wire \sdram|m_addr[12]~q ;
wire \sdram|m_bank[0]~q ;
wire \sdram|m_bank[1]~q ;
wire \sdram|m_cmd[1]~q ;
wire \sdram|m_cmd[3]~q ;
wire \sdram|m_dqm[0]~q ;
wire \sdram|m_dqm[1]~q ;
wire \sdram|m_dqm[2]~q ;
wire \sdram|m_dqm[3]~q ;
wire \sdram|m_cmd[2]~q ;
wire \sdram|m_cmd[0]~q ;
wire \jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|adapted_tdo~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|sr[0]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[0]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[1]~q ;
wire \nios2|cpu|d_writedata[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \nios2|cpu|d_write~q ;
wire \mm_interconnect_0|nios2_data_master_translator|write_accepted~q ;
wire \led|always0~0_combout ;
wire \mm_interconnect_0|router|Equal4~1_combout ;
wire \jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|rst1~q ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ;
wire \led|always0~1_combout ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \nios2|cpu|d_writedata[1]~q ;
wire \nios2|cpu|d_writedata[2]~q ;
wire \nios2|cpu|d_writedata[3]~q ;
wire \nios2|cpu|d_writedata[4]~q ;
wire \nios2|cpu|d_writedata[5]~q ;
wire \nios2|cpu|d_writedata[6]~q ;
wire \nios2|cpu|d_writedata[7]~q ;
wire \sdram|the_sdram_demo_sdram_input_efifo_module|entries[1]~q ;
wire \sdram|the_sdram_demo_sdram_input_efifo_module|entries[0]~q ;
wire \nios2|cpu|d_read~q ;
wire \mm_interconnect_0|nios2_data_master_translator|av_waitrequest~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_begintransfer~0_combout ;
wire \mm_interconnect_0|cmd_demux|sink_ready~1_combout ;
wire \mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_demux|WideOr0~0_combout ;
wire \mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ;
wire \mm_interconnect_0|ram_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal5~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_demux|WideOr0~4_combout ;
wire \mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ;
wire \sdram|za_valid~q ;
wire \mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|nios2_data_master_translator|av_waitrequest~1_combout ;
wire \mm_interconnect_0|router|Equal1~3_combout ;
wire \mm_interconnect_0|cmd_demux|src5_valid~1_combout ;
wire \mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ;
wire \nios2|cpu|i_read~q ;
wire \nios2|cpu|F_pc[25]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[68]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[58]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_valid~1_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[59]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[60]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[61]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[62]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[51]~combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~0_combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~1_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[52]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[53]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[54]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[55]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[56]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[57]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[47]~combout ;
wire \nios2|cpu|d_byteenable[0]~q ;
wire \nios2|cpu|d_byteenable[1]~q ;
wire \nios2|cpu|d_byteenable[2]~q ;
wire \nios2|cpu|d_byteenable[3]~q ;
wire \sdram|m_data[0]~q ;
wire \sdram|m_data[1]~q ;
wire \sdram|m_data[2]~q ;
wire \sdram|m_data[3]~q ;
wire \sdram|m_data[4]~q ;
wire \sdram|m_data[5]~q ;
wire \sdram|m_data[6]~q ;
wire \sdram|m_data[7]~q ;
wire \sdram|m_data[8]~q ;
wire \sdram|m_data[9]~q ;
wire \sdram|m_data[10]~q ;
wire \sdram|m_data[11]~q ;
wire \sdram|m_data[12]~q ;
wire \sdram|m_data[13]~q ;
wire \sdram|m_data[14]~q ;
wire \sdram|m_data[15]~q ;
wire \sdram|m_data[16]~q ;
wire \sdram|m_data[17]~q ;
wire \sdram|m_data[18]~q ;
wire \sdram|m_data[19]~q ;
wire \sdram|m_data[20]~q ;
wire \sdram|m_data[21]~q ;
wire \sdram|m_data[22]~q ;
wire \sdram|m_data[23]~q ;
wire \sdram|m_data[24]~q ;
wire \sdram|m_data[25]~q ;
wire \sdram|m_data[26]~q ;
wire \sdram|m_data[27]~q ;
wire \sdram|m_data[28]~q ;
wire \sdram|m_data[29]~q ;
wire \sdram|m_data[30]~q ;
wire \sdram|m_data[31]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_valid~0_combout ;
wire \mm_interconnect_0|nios2_debug_mem_slave_agent|rf_source_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ;
wire \nios2|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \sdram|za_data[0]~q ;
wire \ram|the_altsyncram|auto_generated|address_reg_a[0]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~1_combout ;
wire \sdram|za_data[22]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \sdram|za_data[23]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \sdram|za_data[24]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \sdram|za_data[25]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \sdram|za_data[26]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \sdram|za_data[1]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \sdram|za_data[4]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \sdram|za_data[3]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \sdram|za_data[2]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[46]~combout ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \sdram|za_data[11]~q ;
wire \sdram|za_data[12]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \sdram|za_data[13]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \sdram|za_data[14]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \sdram|za_data[15]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \sdram|za_data[16]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \sdram|za_data[5]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \sdram|za_data[8]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \sdram|za_data[10]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \sdram|za_data[9]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \sdram|za_data[28]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \sdram|za_data[21]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \sdram|za_data[29]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \sdram|za_data[30]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \sdram|za_data[31]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \sdram|za_data[17]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \sdram|za_data[18]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \sdram|za_data[27]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \sdram|za_data[7]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \sdram|za_data[6]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \sdram|za_data[20]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \sdram|za_data[19]~q ;
wire \mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~3_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~5_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~7_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~9_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~11_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~13_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~15_combout ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~23_combout ;
wire \nios2|cpu|d_writedata[24]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~24_combout ;
wire \nios2|cpu|d_writedata[25]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~25_combout ;
wire \nios2|cpu|d_writedata[26]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~26_combout ;
wire \nios2|cpu|d_writedata[27]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~27_combout ;
wire \nios2|cpu|d_writedata[28]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~28_combout ;
wire \nios2|cpu|d_writedata[29]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~29_combout ;
wire \nios2|cpu|d_writedata[30]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~30_combout ;
wire \nios2|cpu|d_writedata[31]~q ;
wire \mm_interconnect_0|cmd_mux_005|src_payload~31_combout ;
wire \sw|readdata[0]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_data[51]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[32]~combout ;
wire \jtag_uart|ien_AF~q ;
wire \jtag_uart|read_0~q ;
wire \led|readdata[0]~combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \jtag_uart|ien_AE~q ;
wire \jtag_uart|av_readdata[9]~combout ;
wire \jtag_uart|av_readdata[8]~0_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~19_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~20_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[24]~16_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~22_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[25]~17_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~23_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[26]~18_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~24_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[27]~19_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~25_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[28]~20_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~30_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~31_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \sw|readdata[1]~q ;
wire \led|readdata[1]~combout ;
wire \sw|readdata[2]~q ;
wire \led|readdata[2]~combout ;
wire \sw|readdata[3]~q ;
wire \led|readdata[3]~combout ;
wire \sw|readdata[4]~q ;
wire \led|readdata[4]~combout ;
wire \sw|readdata[5]~q ;
wire \led|readdata[5]~combout ;
wire \sw|readdata[6]~q ;
wire \led|readdata[6]~combout ;
wire \sw|readdata[7]~q ;
wire \led|readdata[7]~combout ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[32]~combout ;
wire \jtag_uart|the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \mm_interconnect_0|rsp_mux|src_data[29]~21_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[30]~22_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[31]~23_combout ;
wire \jtag_uart|rvalid~q ;
wire \jtag_uart|woverflow~q ;
wire \jtag_uart|ac~q ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~3_combout ;
wire \nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|resetrequest~q ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \sdram_wire_dq[0]~input_o ;
wire \sdram_wire_dq[1]~input_o ;
wire \sdram_wire_dq[2]~input_o ;
wire \sdram_wire_dq[3]~input_o ;
wire \sdram_wire_dq[4]~input_o ;
wire \sdram_wire_dq[5]~input_o ;
wire \sdram_wire_dq[6]~input_o ;
wire \sdram_wire_dq[7]~input_o ;
wire \sdram_wire_dq[8]~input_o ;
wire \sdram_wire_dq[9]~input_o ;
wire \sdram_wire_dq[10]~input_o ;
wire \sdram_wire_dq[11]~input_o ;
wire \sdram_wire_dq[12]~input_o ;
wire \sdram_wire_dq[13]~input_o ;
wire \sdram_wire_dq[14]~input_o ;
wire \sdram_wire_dq[15]~input_o ;
wire \sdram_wire_dq[16]~input_o ;
wire \sdram_wire_dq[17]~input_o ;
wire \sdram_wire_dq[18]~input_o ;
wire \sdram_wire_dq[19]~input_o ;
wire \sdram_wire_dq[20]~input_o ;
wire \sdram_wire_dq[21]~input_o ;
wire \sdram_wire_dq[22]~input_o ;
wire \sdram_wire_dq[23]~input_o ;
wire \sdram_wire_dq[24]~input_o ;
wire \sdram_wire_dq[25]~input_o ;
wire \sdram_wire_dq[26]~input_o ;
wire \sdram_wire_dq[27]~input_o ;
wire \sdram_wire_dq[28]~input_o ;
wire \sdram_wire_dq[29]~input_o ;
wire \sdram_wire_dq[30]~input_o ;
wire \sdram_wire_dq[31]~input_o ;
wire \clk_clk~input_o ;
wire \sw_export[0]~input_o ;
wire \sw_export[1]~input_o ;
wire \sw_export[2]~input_o ;
wire \sw_export[3]~input_o ;
wire \sw_export[4]~input_o ;
wire \sw_export[5]~input_o ;
wire \sw_export[6]~input_o ;
wire \sw_export[7]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


sdram_demo_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.resetrequest(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|resetrequest~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_jtag_uart jtag_uart(
	.W_alu_result_2(\nios2|cpu|W_alu_result[2]~q ),
	.d_writedata_10(\nios2|cpu|d_writedata[10]~q ),
	.q_b_0(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.adapted_tdo(\jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|adapted_tdo~q ),
	.d_writedata_0(\nios2|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.always0(\led|always0~0_combout ),
	.rst1(\jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|rst1~q ),
	.d_writedata_1(\nios2|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2|cpu|d_writedata[7]~q ),
	.av_begintransfer(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_begintransfer~0_combout ),
	.Equal5(\mm_interconnect_0|router|Equal5~1_combout ),
	.av_waitrequest1(\jtag_uart|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.b_full(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.ien_AF1(\jtag_uart|ien_AF~q ),
	.read_01(\jtag_uart|read_0~q ),
	.ien_AE1(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.b_non_empty(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.b_full1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.rvalid1(\jtag_uart|rvalid~q ),
	.woverflow1(\jtag_uart|woverflow~q ),
	.ac1(\jtag_uart|ac~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_nios2 nios2(
	.W_alu_result_4(\nios2|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\nios2|cpu|W_alu_result[5]~q ),
	.W_alu_result_9(\nios2|cpu|W_alu_result[9]~q ),
	.W_alu_result_24(\nios2|cpu|W_alu_result[24]~q ),
	.W_alu_result_25(\nios2|cpu|W_alu_result[25]~q ),
	.W_alu_result_26(\nios2|cpu|W_alu_result[26]~q ),
	.W_alu_result_27(\nios2|cpu|W_alu_result[27]~q ),
	.W_alu_result_28(\nios2|cpu|W_alu_result[28]~q ),
	.W_alu_result_20(\nios2|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\nios2|cpu|W_alu_result[19]~q ),
	.W_alu_result_21(\nios2|cpu|W_alu_result[21]~q ),
	.W_alu_result_22(\nios2|cpu|W_alu_result[22]~q ),
	.W_alu_result_23(\nios2|cpu|W_alu_result[23]~q ),
	.W_alu_result_18(\nios2|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\nios2|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\nios2|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2|cpu|W_alu_result[13]~q ),
	.W_alu_result_6(\nios2|cpu|W_alu_result[6]~q ),
	.W_alu_result_7(\nios2|cpu|W_alu_result[7]~q ),
	.W_alu_result_8(\nios2|cpu|W_alu_result[8]~q ),
	.W_alu_result_12(\nios2|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\nios2|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2|cpu|W_alu_result[10]~q ),
	.W_alu_result_2(\nios2|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2|cpu|W_alu_result[3]~q ),
	.F_pc_17(\nios2|cpu|F_pc[17]~q ),
	.F_pc_16(\nios2|cpu|F_pc[16]~q ),
	.F_pc_18(\nios2|cpu|F_pc[18]~q ),
	.F_pc_19(\nios2|cpu|F_pc[19]~q ),
	.F_pc_20(\nios2|cpu|F_pc[20]~q ),
	.F_pc_21(\nios2|cpu|F_pc[21]~q ),
	.F_pc_22(\nios2|cpu|F_pc[22]~q ),
	.F_pc_23(\nios2|cpu|F_pc[23]~q ),
	.F_pc_24(\nios2|cpu|F_pc[24]~q ),
	.F_pc_26(\nios2|cpu|F_pc[26]~q ),
	.F_pc_15(\nios2|cpu|F_pc[15]~q ),
	.F_pc_14(\nios2|cpu|F_pc[14]~q ),
	.F_pc_9(\nios2|cpu|F_pc[9]~q ),
	.F_pc_11(\nios2|cpu|F_pc[11]~q ),
	.F_pc_13(\nios2|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2|cpu|F_pc[12]~q ),
	.F_pc_10(\nios2|cpu|F_pc[10]~q ),
	.F_pc_0(\nios2|cpu|F_pc[0]~q ),
	.F_pc_1(\nios2|cpu|F_pc[1]~q ),
	.F_pc_2(\nios2|cpu|F_pc[2]~q ),
	.F_pc_3(\nios2|cpu|F_pc[3]~q ),
	.F_pc_4(\nios2|cpu|F_pc[4]~q ),
	.F_pc_5(\nios2|cpu|F_pc[5]~q ),
	.F_pc_6(\nios2|cpu|F_pc[6]~q ),
	.F_pc_7(\nios2|cpu|F_pc[7]~q ),
	.F_pc_8(\nios2|cpu|F_pc[8]~q ),
	.ram_block1a32(\ram|the_altsyncram|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a0(\ram|the_altsyncram|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a54(\ram|the_altsyncram|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a22(\ram|the_altsyncram|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a55(\ram|the_altsyncram|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a23(\ram|the_altsyncram|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a56(\ram|the_altsyncram|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a24(\ram|the_altsyncram|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a57(\ram|the_altsyncram|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a25(\ram|the_altsyncram|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a58(\ram|the_altsyncram|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a26(\ram|the_altsyncram|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a33(\ram|the_altsyncram|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a1(\ram|the_altsyncram|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a36(\ram|the_altsyncram|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a4(\ram|the_altsyncram|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a35(\ram|the_altsyncram|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a3(\ram|the_altsyncram|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a34(\ram|the_altsyncram|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a2(\ram|the_altsyncram|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a43(\ram|the_altsyncram|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a11(\ram|the_altsyncram|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a44(\ram|the_altsyncram|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a12(\ram|the_altsyncram|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a45(\ram|the_altsyncram|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a13(\ram|the_altsyncram|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a46(\ram|the_altsyncram|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a14(\ram|the_altsyncram|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a47(\ram|the_altsyncram|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a15(\ram|the_altsyncram|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a48(\ram|the_altsyncram|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a16(\ram|the_altsyncram|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a37(\ram|the_altsyncram|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a5(\ram|the_altsyncram|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a40(\ram|the_altsyncram|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a8(\ram|the_altsyncram|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a42(\ram|the_altsyncram|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a10(\ram|the_altsyncram|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a41(\ram|the_altsyncram|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a9(\ram|the_altsyncram|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a60(\ram|the_altsyncram|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a28(\ram|the_altsyncram|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a53(\ram|the_altsyncram|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a21(\ram|the_altsyncram|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a61(\ram|the_altsyncram|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a29(\ram|the_altsyncram|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a62(\ram|the_altsyncram|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a30(\ram|the_altsyncram|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a63(\ram|the_altsyncram|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a31(\ram|the_altsyncram|auto_generated|ram_block1a31~portadataout ),
	.ram_block1a49(\ram|the_altsyncram|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a17(\ram|the_altsyncram|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a50(\ram|the_altsyncram|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a18(\ram|the_altsyncram|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a59(\ram|the_altsyncram|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a27(\ram|the_altsyncram|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a39(\ram|the_altsyncram|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a7(\ram|the_altsyncram|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a38(\ram|the_altsyncram|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a6(\ram|the_altsyncram|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a52(\ram|the_altsyncram|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a20(\ram|the_altsyncram|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a51(\ram|the_altsyncram|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a19(\ram|the_altsyncram|auto_generated|ram_block1a19~portadataout ),
	.d_writedata_8(\nios2|cpu|d_writedata[8]~q ),
	.d_writedata_9(\nios2|cpu|d_writedata[9]~q ),
	.d_writedata_10(\nios2|cpu|d_writedata[10]~q ),
	.d_writedata_11(\nios2|cpu|d_writedata[11]~q ),
	.d_writedata_12(\nios2|cpu|d_writedata[12]~q ),
	.d_writedata_13(\nios2|cpu|d_writedata[13]~q ),
	.d_writedata_14(\nios2|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios2|cpu|d_writedata[15]~q ),
	.d_writedata_16(\nios2|cpu|d_writedata[16]~q ),
	.d_writedata_17(\nios2|cpu|d_writedata[17]~q ),
	.d_writedata_18(\nios2|cpu|d_writedata[18]~q ),
	.d_writedata_19(\nios2|cpu|d_writedata[19]~q ),
	.d_writedata_20(\nios2|cpu|d_writedata[20]~q ),
	.d_writedata_21(\nios2|cpu|d_writedata[21]~q ),
	.d_writedata_22(\nios2|cpu|d_writedata[22]~q ),
	.d_writedata_23(\nios2|cpu|d_writedata[23]~q ),
	.readdata_0(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[0]~q ),
	.readdata_22(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[23]~q ),
	.readdata_24(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[26]~q ),
	.readdata_1(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[1]~q ),
	.readdata_4(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[4]~q ),
	.readdata_3(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[2]~q ),
	.readdata_11(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[11]~q ),
	.readdata_12(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[12]~q ),
	.readdata_13(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[13]~q ),
	.readdata_14(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[15]~q ),
	.readdata_16(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[16]~q ),
	.readdata_5(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[5]~q ),
	.readdata_8(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[8]~q ),
	.readdata_10(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[10]~q ),
	.readdata_9(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[9]~q ),
	.readdata_28(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[28]~q ),
	.readdata_21(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[21]~q ),
	.readdata_29(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[31]~q ),
	.readdata_17(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[17]~q ),
	.readdata_18(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[18]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.readdata_27(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[27]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.readdata_7(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[6]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.readdata_20(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[20]~q ),
	.readdata_19(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[19]~q ),
	.sr_0(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|sr[0]~q ),
	.ir_out_0(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_writedata_0(\nios2|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_write(\nios2|cpu|d_write~q ),
	.always0(\led|always0~0_combout ),
	.d_writedata_1(\nios2|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2|cpu|d_writedata[7]~q ),
	.d_read(\nios2|cpu|d_read~q ),
	.av_waitrequest(\mm_interconnect_0|nios2_data_master_translator|av_waitrequest~0_combout ),
	.sink_ready(\mm_interconnect_0|cmd_demux|sink_ready~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~4_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.av_waitrequest1(\mm_interconnect_0|nios2_data_master_translator|av_waitrequest~1_combout ),
	.i_read(\nios2|cpu|i_read~q ),
	.F_pc_25(\nios2|cpu|F_pc[25]~q ),
	.d_byteenable_0(\nios2|cpu|d_byteenable[0]~q ),
	.d_byteenable_1(\nios2|cpu|d_byteenable[1]~q ),
	.d_byteenable_2(\nios2|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\nios2|cpu|d_byteenable[3]~q ),
	.rf_source_valid(\mm_interconnect_0|nios2_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.hbreak_enabled(\nios2|cpu|hbreak_enabled~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.address_reg_a_0(\ram|the_altsyncram|auto_generated|address_reg_a[0]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~1_combout ),
	.za_data_22(\sdram|za_data[22]~q ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.WideOr13(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~3_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~5_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~7_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~9_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~11_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~13_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~15_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.d_writedata_24(\nios2|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios2|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios2|cpu|d_writedata[26]~q ),
	.d_writedata_27(\nios2|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios2|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios2|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios2|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios2|cpu|d_writedata[31]~q ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.src_data_24(\mm_interconnect_0|rsp_mux|src_data[24]~16_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux|src_data[25]~17_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux|src_data[26]~18_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux|src_data[27]~19_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux|src_data[28]~20_combout ),
	.av_readdata_pre_151(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_141(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_131(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_121(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux|src_data[29]~21_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux|src_data[30]~22_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[31]~23_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.debug_reset_request(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|resetrequest~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_led led(
	.W_alu_result_4(\nios2|cpu|W_alu_result[4]~q ),
	.W_alu_result_2(\nios2|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2|cpu|W_alu_result[3]~q ),
	.data_out_0(\led|data_out[0]~q ),
	.data_out_1(\led|data_out[1]~q ),
	.data_out_2(\led|data_out[2]~q ),
	.data_out_3(\led|data_out[3]~q ),
	.data_out_4(\led|data_out[4]~q ),
	.data_out_5(\led|data_out[5]~q ),
	.data_out_6(\led|data_out[6]~q ),
	.data_out_7(\led|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2|cpu|d_writedata[7]~q ,\nios2|cpu|d_writedata[6]~q ,\nios2|cpu|d_writedata[5]~q ,\nios2|cpu|d_writedata[4]~q ,\nios2|cpu|d_writedata[3]~q ,\nios2|cpu|d_writedata[2]~q ,
\nios2|cpu|d_writedata[1]~q ,\nios2|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.d_write(\nios2|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_data_master_translator|write_accepted~q ),
	.always0(\led|always0~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~1_combout ),
	.rst1(\jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|rst1~q ),
	.wait_latency_counter_1(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.always01(\led|always0~1_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.mem_used_1(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.readdata_0(\led|readdata[0]~combout ),
	.readdata_1(\led|readdata[1]~combout ),
	.readdata_2(\led|readdata[2]~combout ),
	.readdata_3(\led|readdata[3]~combout ),
	.readdata_4(\led|readdata[4]~combout ),
	.readdata_5(\led|readdata[5]~combout ),
	.readdata_6(\led|readdata[6]~combout ),
	.readdata_7(\led|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_ram ram(
	.ram_block1a32(\ram|the_altsyncram|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a0(\ram|the_altsyncram|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a54(\ram|the_altsyncram|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a22(\ram|the_altsyncram|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a55(\ram|the_altsyncram|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a23(\ram|the_altsyncram|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a56(\ram|the_altsyncram|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a24(\ram|the_altsyncram|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a57(\ram|the_altsyncram|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a25(\ram|the_altsyncram|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a58(\ram|the_altsyncram|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a26(\ram|the_altsyncram|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a33(\ram|the_altsyncram|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a1(\ram|the_altsyncram|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a36(\ram|the_altsyncram|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a4(\ram|the_altsyncram|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a35(\ram|the_altsyncram|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a3(\ram|the_altsyncram|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a34(\ram|the_altsyncram|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a2(\ram|the_altsyncram|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a43(\ram|the_altsyncram|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a11(\ram|the_altsyncram|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a44(\ram|the_altsyncram|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a12(\ram|the_altsyncram|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a45(\ram|the_altsyncram|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a13(\ram|the_altsyncram|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a46(\ram|the_altsyncram|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a14(\ram|the_altsyncram|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a47(\ram|the_altsyncram|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a15(\ram|the_altsyncram|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a48(\ram|the_altsyncram|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a16(\ram|the_altsyncram|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a37(\ram|the_altsyncram|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a5(\ram|the_altsyncram|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a40(\ram|the_altsyncram|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a8(\ram|the_altsyncram|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a42(\ram|the_altsyncram|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a10(\ram|the_altsyncram|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a41(\ram|the_altsyncram|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a9(\ram|the_altsyncram|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a60(\ram|the_altsyncram|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a28(\ram|the_altsyncram|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a53(\ram|the_altsyncram|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a21(\ram|the_altsyncram|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a61(\ram|the_altsyncram|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a29(\ram|the_altsyncram|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a62(\ram|the_altsyncram|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a30(\ram|the_altsyncram|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a63(\ram|the_altsyncram|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a31(\ram|the_altsyncram|auto_generated|ram_block1a31~portadataout ),
	.ram_block1a49(\ram|the_altsyncram|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a17(\ram|the_altsyncram|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a50(\ram|the_altsyncram|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a18(\ram|the_altsyncram|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a59(\ram|the_altsyncram|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a27(\ram|the_altsyncram|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a39(\ram|the_altsyncram|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a7(\ram|the_altsyncram|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a38(\ram|the_altsyncram|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a6(\ram|the_altsyncram|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a52(\ram|the_altsyncram|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a20(\ram|the_altsyncram|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a51(\ram|the_altsyncram|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a19(\ram|the_altsyncram|auto_generated|ram_block1a19~portadataout ),
	.d_write(\nios2|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_data_master_translator|write_accepted~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~3_combout ),
	.src5_valid(\mm_interconnect_0|cmd_demux|src5_valid~1_combout ),
	.src_valid(\mm_interconnect_0|cmd_mux_004|src_valid~0_combout ),
	.address_reg_a_0(\ram|the_altsyncram|auto_generated|address_reg_a[0]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_data_51(\mm_interconnect_0|cmd_mux_004|src_data[51]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_004|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_004|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_004|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_004|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_004|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_004|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_004|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_004|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_004|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_004|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_004|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_004|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_004|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_004|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_004|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_004|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_004|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_004|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_004|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_004|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_004|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_004|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_004|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_004|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_004|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_004|src_payload~10_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_004|src_data[33]~combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_004|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_004|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_004|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_004|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_004|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_004|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_004|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_004|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_004|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_004|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_004|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_004|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_004|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_004|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_004|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_004|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_004|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_004|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_004|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_004|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_004|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_mm_interconnect_0 mm_interconnect_0(
	.W_alu_result_4(\nios2|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\nios2|cpu|W_alu_result[5]~q ),
	.W_alu_result_9(\nios2|cpu|W_alu_result[9]~q ),
	.W_alu_result_24(\nios2|cpu|W_alu_result[24]~q ),
	.W_alu_result_25(\nios2|cpu|W_alu_result[25]~q ),
	.W_alu_result_26(\nios2|cpu|W_alu_result[26]~q ),
	.W_alu_result_27(\nios2|cpu|W_alu_result[27]~q ),
	.W_alu_result_28(\nios2|cpu|W_alu_result[28]~q ),
	.W_alu_result_20(\nios2|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\nios2|cpu|W_alu_result[19]~q ),
	.W_alu_result_21(\nios2|cpu|W_alu_result[21]~q ),
	.W_alu_result_22(\nios2|cpu|W_alu_result[22]~q ),
	.W_alu_result_23(\nios2|cpu|W_alu_result[23]~q ),
	.W_alu_result_18(\nios2|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\nios2|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\nios2|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2|cpu|W_alu_result[13]~q ),
	.W_alu_result_6(\nios2|cpu|W_alu_result[6]~q ),
	.W_alu_result_7(\nios2|cpu|W_alu_result[7]~q ),
	.W_alu_result_8(\nios2|cpu|W_alu_result[8]~q ),
	.W_alu_result_12(\nios2|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\nios2|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2|cpu|W_alu_result[10]~q ),
	.W_alu_result_2(\nios2|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2|cpu|W_alu_result[3]~q ),
	.F_pc_17(\nios2|cpu|F_pc[17]~q ),
	.F_pc_16(\nios2|cpu|F_pc[16]~q ),
	.F_pc_18(\nios2|cpu|F_pc[18]~q ),
	.F_pc_19(\nios2|cpu|F_pc[19]~q ),
	.F_pc_20(\nios2|cpu|F_pc[20]~q ),
	.F_pc_21(\nios2|cpu|F_pc[21]~q ),
	.F_pc_22(\nios2|cpu|F_pc[22]~q ),
	.F_pc_23(\nios2|cpu|F_pc[23]~q ),
	.F_pc_24(\nios2|cpu|F_pc[24]~q ),
	.F_pc_26(\nios2|cpu|F_pc[26]~q ),
	.F_pc_15(\nios2|cpu|F_pc[15]~q ),
	.F_pc_14(\nios2|cpu|F_pc[14]~q ),
	.F_pc_9(\nios2|cpu|F_pc[9]~q ),
	.F_pc_11(\nios2|cpu|F_pc[11]~q ),
	.F_pc_13(\nios2|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2|cpu|F_pc[12]~q ),
	.F_pc_10(\nios2|cpu|F_pc[10]~q ),
	.F_pc_0(\nios2|cpu|F_pc[0]~q ),
	.F_pc_1(\nios2|cpu|F_pc[1]~q ),
	.F_pc_2(\nios2|cpu|F_pc[2]~q ),
	.F_pc_3(\nios2|cpu|F_pc[3]~q ),
	.F_pc_4(\nios2|cpu|F_pc[4]~q ),
	.F_pc_5(\nios2|cpu|F_pc[5]~q ),
	.F_pc_6(\nios2|cpu|F_pc[6]~q ),
	.F_pc_7(\nios2|cpu|F_pc[7]~q ),
	.F_pc_8(\nios2|cpu|F_pc[8]~q ),
	.ram_block1a32(\ram|the_altsyncram|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a0(\ram|the_altsyncram|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a56(\ram|the_altsyncram|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a24(\ram|the_altsyncram|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a57(\ram|the_altsyncram|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a25(\ram|the_altsyncram|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a58(\ram|the_altsyncram|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a26(\ram|the_altsyncram|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a33(\ram|the_altsyncram|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a1(\ram|the_altsyncram|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a36(\ram|the_altsyncram|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a4(\ram|the_altsyncram|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a35(\ram|the_altsyncram|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a3(\ram|the_altsyncram|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a34(\ram|the_altsyncram|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a2(\ram|the_altsyncram|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a37(\ram|the_altsyncram|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a5(\ram|the_altsyncram|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a60(\ram|the_altsyncram|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a28(\ram|the_altsyncram|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a61(\ram|the_altsyncram|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a29(\ram|the_altsyncram|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a62(\ram|the_altsyncram|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a30(\ram|the_altsyncram|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a63(\ram|the_altsyncram|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a31(\ram|the_altsyncram|auto_generated|ram_block1a31~portadataout ),
	.ram_block1a59(\ram|the_altsyncram|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a27(\ram|the_altsyncram|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a39(\ram|the_altsyncram|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a7(\ram|the_altsyncram|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a38(\ram|the_altsyncram|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a6(\ram|the_altsyncram|auto_generated|ram_block1a6~portadataout ),
	.d_writedata_8(\nios2|cpu|d_writedata[8]~q ),
	.d_writedata_9(\nios2|cpu|d_writedata[9]~q ),
	.d_writedata_10(\nios2|cpu|d_writedata[10]~q ),
	.d_writedata_11(\nios2|cpu|d_writedata[11]~q ),
	.d_writedata_12(\nios2|cpu|d_writedata[12]~q ),
	.d_writedata_13(\nios2|cpu|d_writedata[13]~q ),
	.d_writedata_14(\nios2|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios2|cpu|d_writedata[15]~q ),
	.d_writedata_16(\nios2|cpu|d_writedata[16]~q ),
	.d_writedata_17(\nios2|cpu|d_writedata[17]~q ),
	.d_writedata_18(\nios2|cpu|d_writedata[18]~q ),
	.d_writedata_19(\nios2|cpu|d_writedata[19]~q ),
	.d_writedata_20(\nios2|cpu|d_writedata[20]~q ),
	.d_writedata_21(\nios2|cpu|d_writedata[21]~q ),
	.d_writedata_22(\nios2|cpu|d_writedata[22]~q ),
	.d_writedata_23(\nios2|cpu|d_writedata[23]~q ),
	.readdata_0(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[0]~q ),
	.q_b_0(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.readdata_22(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[23]~q ),
	.readdata_24(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[26]~q ),
	.readdata_1(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[1]~q ),
	.readdata_4(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[4]~q ),
	.readdata_3(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[2]~q ),
	.readdata_11(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[11]~q ),
	.readdata_12(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[12]~q ),
	.readdata_13(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[13]~q ),
	.readdata_14(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[15]~q ),
	.readdata_16(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[16]~q ),
	.readdata_5(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[5]~q ),
	.readdata_8(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[8]~q ),
	.readdata_10(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[10]~q ),
	.readdata_9(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[9]~q ),
	.readdata_28(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[28]~q ),
	.readdata_21(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[21]~q ),
	.readdata_29(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[31]~q ),
	.readdata_17(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[17]~q ),
	.readdata_18(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[18]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.readdata_27(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[27]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.readdata_7(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[6]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.readdata_20(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[20]~q ),
	.readdata_19(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|readdata[19]~q ),
	.q_b_1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.d_writedata_0(\nios2|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_write(\nios2|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_data_master_translator|write_accepted~q ),
	.always0(\led|always0~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~1_combout ),
	.rst1(\jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|rst1~q ),
	.wait_latency_counter_1(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.always01(\led|always0~1_combout ),
	.wait_latency_counter_0(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.mem_used_1(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.d_writedata_1(\nios2|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2|cpu|d_writedata[7]~q ),
	.entries_1(\sdram|the_sdram_demo_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_sdram_demo_sdram_input_efifo_module|entries[0]~q ),
	.d_read(\nios2|cpu|d_read~q ),
	.nios2_data_master_waitrequest(\mm_interconnect_0|nios2_data_master_translator|av_waitrequest~0_combout ),
	.av_begintransfer(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_begintransfer~0_combout ),
	.sink_ready(\mm_interconnect_0|cmd_demux|sink_ready~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~0_combout ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_004|saved_grant[0]~q ),
	.mem_used_11(\mm_interconnect_0|ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal5(\mm_interconnect_0|router|Equal5~1_combout ),
	.saved_grant_02(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.waitrequest(\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_12(\mm_interconnect_0|nios2_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\jtag_uart|av_waitrequest~q ),
	.mem_used_13(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr01(\mm_interconnect_0|cmd_demux|WideOr0~4_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.za_valid(\sdram|za_valid~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.av_waitrequest1(\mm_interconnect_0|nios2_data_master_translator|av_waitrequest~1_combout ),
	.Equal1(\mm_interconnect_0|router|Equal1~3_combout ),
	.src5_valid(\mm_interconnect_0|cmd_demux|src5_valid~1_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ),
	.i_read(\nios2|cpu|i_read~q ),
	.F_pc_25(\nios2|cpu|F_pc[25]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_005|src_valid~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_005|src_data[68]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_005|src_data[58]~combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_005|src_valid~1_combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_005|src_data[59]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_005|src_data[60]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_005|src_data[61]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_005|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_005|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_005|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_005|src_data[50]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_005|src_data[51]~combout ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~0_combout ),
	.m0_write1(\mm_interconnect_0|sdram_s1_agent|m0_write~1_combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_005|src_data[52]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_005|src_data[53]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_005|src_data[54]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_005|src_data[55]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_005|src_data[56]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_005|src_data[57]~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_005|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_005|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_005|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_005|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_005|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_005|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_005|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_005|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_005|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_005|src_data[47]~combout ),
	.d_byteenable_0(\nios2|cpu|d_byteenable[0]~q ),
	.d_byteenable_1(\nios2|cpu|d_byteenable[1]~q ),
	.d_byteenable_2(\nios2|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\nios2|cpu|d_byteenable[3]~q ),
	.src_valid2(\mm_interconnect_0|cmd_mux_004|src_valid~0_combout ),
	.rf_source_valid(\mm_interconnect_0|nios2_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_005|src1_valid~0_combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.hbreak_enabled(\nios2|cpu|hbreak_enabled~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.address_reg_a_0(\ram|the_altsyncram|auto_generated|address_reg_a[0]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~1_combout ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.WideOr13(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~3_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~5_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~7_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~9_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~11_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~13_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~15_combout ),
	.b_full(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_005|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_005|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_005|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_005|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_005|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_005|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_005|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_005|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_005|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_005|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_005|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_005|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_005|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_005|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_005|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_005|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_005|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_005|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_005|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_005|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_005|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_005|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_005|src_payload~23_combout ),
	.d_writedata_24(\nios2|cpu|d_writedata[24]~q ),
	.src_payload24(\mm_interconnect_0|cmd_mux_005|src_payload~24_combout ),
	.d_writedata_25(\nios2|cpu|d_writedata[25]~q ),
	.src_payload25(\mm_interconnect_0|cmd_mux_005|src_payload~25_combout ),
	.d_writedata_26(\nios2|cpu|d_writedata[26]~q ),
	.src_payload26(\mm_interconnect_0|cmd_mux_005|src_payload~26_combout ),
	.d_writedata_27(\nios2|cpu|d_writedata[27]~q ),
	.src_payload27(\mm_interconnect_0|cmd_mux_005|src_payload~27_combout ),
	.d_writedata_28(\nios2|cpu|d_writedata[28]~q ),
	.src_payload28(\mm_interconnect_0|cmd_mux_005|src_payload~28_combout ),
	.d_writedata_29(\nios2|cpu|d_writedata[29]~q ),
	.src_payload29(\mm_interconnect_0|cmd_mux_005|src_payload~29_combout ),
	.d_writedata_30(\nios2|cpu|d_writedata[30]~q ),
	.src_payload30(\mm_interconnect_0|cmd_mux_005|src_payload~30_combout ),
	.d_writedata_31(\nios2|cpu|d_writedata[31]~q ),
	.src_payload31(\mm_interconnect_0|cmd_mux_005|src_payload~31_combout ),
	.readdata_01(\sw|readdata[0]~q ),
	.src_data_511(\mm_interconnect_0|cmd_mux_004|src_data[51]~combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_004|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_004|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_004|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_004|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_004|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_004|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_004|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_004|src_data[45]~combout ),
	.src_data_462(\mm_interconnect_0|cmd_mux_004|src_data[46]~combout ),
	.src_data_471(\mm_interconnect_0|cmd_mux_004|src_data[47]~combout ),
	.src_data_481(\mm_interconnect_0|cmd_mux_004|src_data[48]~combout ),
	.src_data_491(\mm_interconnect_0|cmd_mux_004|src_data[49]~combout ),
	.src_data_501(\mm_interconnect_0|cmd_mux_004|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_004|src_data[32]~combout ),
	.ien_AF(\jtag_uart|ien_AF~q ),
	.read_0(\jtag_uart|read_0~q ),
	.readdata_02(\led|readdata[0]~combout ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.ien_AE(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_004|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_004|src_data[34]~combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_004|src_payload~2_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_004|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_004|src_data[35]~combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_004|src_payload~4_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_004|src_payload~5_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_004|src_payload~6_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_004|src_payload~7_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_004|src_payload~8_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_004|src_payload~9_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_004|src_payload~10_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_004|src_data[33]~combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_004|src_payload~11_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_004|src_payload~12_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_004|src_payload~13_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_004|src_payload~14_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_004|src_payload~15_combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_004|src_payload~16_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_004|src_payload~17_combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_004|src_payload~18_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_004|src_payload~19_combout ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_004|src_payload~20_combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux|src_data[24]~16_combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_004|src_payload~21_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_004|src_payload~22_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux|src_data[25]~17_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_004|src_payload~23_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux|src_data[26]~18_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_004|src_payload~24_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux|src_data[27]~19_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_004|src_payload~25_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux|src_data[28]~20_combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_004|src_payload~26_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_004|src_payload~27_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_004|src_payload~28_combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_004|src_payload~29_combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_004|src_payload~30_combout ),
	.av_readdata_pre_151(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.src_payload63(\mm_interconnect_0|cmd_mux_004|src_payload~31_combout ),
	.av_readdata_pre_141(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_131(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_121(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.readdata_110(\sw|readdata[1]~q ),
	.readdata_111(\led|readdata[1]~combout ),
	.readdata_210(\sw|readdata[2]~q ),
	.readdata_211(\led|readdata[2]~combout ),
	.readdata_32(\sw|readdata[3]~q ),
	.readdata_33(\led|readdata[3]~combout ),
	.readdata_41(\sw|readdata[4]~q ),
	.readdata_42(\led|readdata[4]~combout ),
	.readdata_51(\sw|readdata[5]~q ),
	.readdata_52(\led|readdata[5]~combout ),
	.readdata_61(\sw|readdata[6]~q ),
	.readdata_62(\led|readdata[6]~combout ),
	.readdata_71(\sw|readdata[7]~q ),
	.readdata_72(\led|readdata[7]~combout ),
	.b_non_empty(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.src_payload64(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_data_382(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_402(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_392(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_data_452(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_442(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_432(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_422(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_412(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.b_full1(\jtag_uart|the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_data_29(\mm_interconnect_0|rsp_mux|src_data[29]~21_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux|src_data[30]~22_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[31]~23_combout ),
	.rvalid(\jtag_uart|rvalid~q ),
	.woverflow(\jtag_uart|woverflow~q ),
	.ac(\jtag_uart|ac~q ),
	.src_payload66(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload75(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload76(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload79(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload82(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload83(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload87(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload88(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload89(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload90(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload91(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload92(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload93(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload94(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload95(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload96(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

sdram_demo_sdram_demo_sw sw(
	.W_alu_result_2(\nios2|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2|cpu|W_alu_result[3]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.readdata_0(\sw|readdata[0]~q ),
	.readdata_1(\sw|readdata[1]~q ),
	.readdata_2(\sw|readdata[2]~q ),
	.readdata_3(\sw|readdata[3]~q ),
	.readdata_4(\sw|readdata[4]~q ),
	.readdata_5(\sw|readdata[5]~q ),
	.readdata_6(\sw|readdata[6]~q ),
	.readdata_7(\sw|readdata[7]~q ),
	.clk_clk(\clk_clk~input_o ),
	.sw_export_0(\sw_export[0]~input_o ),
	.sw_export_1(\sw_export[1]~input_o ),
	.sw_export_2(\sw_export[2]~input_o ),
	.sw_export_3(\sw_export[3]~input_o ),
	.sw_export_4(\sw_export[4]~input_o ),
	.sw_export_5(\sw_export[5]~input_o ),
	.sw_export_6(\sw_export[6]~input_o ),
	.sw_export_7(\sw_export[7]~input_o ));

sdram_demo_sdram_demo_sdram sdram(
	.m_addr_0(\sdram|m_addr[0]~q ),
	.m_addr_1(\sdram|m_addr[1]~q ),
	.m_addr_2(\sdram|m_addr[2]~q ),
	.m_addr_3(\sdram|m_addr[3]~q ),
	.m_addr_6(\sdram|m_addr[6]~q ),
	.m_addr_7(\sdram|m_addr[7]~q ),
	.m_addr_8(\sdram|m_addr[8]~q ),
	.m_addr_9(\sdram|m_addr[9]~q ),
	.oe1(\sdram|oe~q ),
	.m_addr_4(\sdram|m_addr[4]~q ),
	.m_addr_5(\sdram|m_addr[5]~q ),
	.m_addr_10(\sdram|m_addr[10]~q ),
	.m_addr_11(\sdram|m_addr[11]~q ),
	.m_addr_12(\sdram|m_addr[12]~q ),
	.m_bank_0(\sdram|m_bank[0]~q ),
	.m_bank_1(\sdram|m_bank[1]~q ),
	.m_cmd_1(\sdram|m_cmd[1]~q ),
	.m_cmd_3(\sdram|m_cmd[3]~q ),
	.m_dqm_0(\sdram|m_dqm[0]~q ),
	.m_dqm_1(\sdram|m_dqm[1]~q ),
	.m_dqm_2(\sdram|m_dqm[2]~q ),
	.m_dqm_3(\sdram|m_dqm[3]~q ),
	.m_cmd_2(\sdram|m_cmd[2]~q ),
	.m_cmd_0(\sdram|m_cmd[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.always0(\led|always0~0_combout ),
	.entries_1(\sdram|the_sdram_demo_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_sdram_demo_sdram_input_efifo_module|entries[0]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_005|saved_grant[0]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~0_combout ),
	.za_valid1(\sdram|za_valid~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~3_combout ),
	.src5_valid(\mm_interconnect_0|cmd_demux|src5_valid~1_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_005|saved_grant[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_005|src_valid~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_005|src_data[68]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_005|src_data[58]~combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_005|src_valid~1_combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_005|src_data[59]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_005|src_data[60]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_005|src_data[61]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_005|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_005|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_005|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_005|src_data[50]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_005|src_data[51]~combout ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~0_combout ),
	.m0_write1(\mm_interconnect_0|sdram_s1_agent|m0_write~1_combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_005|src_data[52]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_005|src_data[53]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_005|src_data[54]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_005|src_data[55]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_005|src_data[56]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_005|src_data[57]~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_005|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_005|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_005|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_005|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_005|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_005|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_005|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_005|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_005|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_005|src_data[47]~combout ),
	.d_byteenable_0(\nios2|cpu|d_byteenable[0]~q ),
	.d_byteenable_1(\nios2|cpu|d_byteenable[1]~q ),
	.d_byteenable_2(\nios2|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\nios2|cpu|d_byteenable[3]~q ),
	.m_data_0(\sdram|m_data[0]~q ),
	.m_data_1(\sdram|m_data[1]~q ),
	.m_data_2(\sdram|m_data[2]~q ),
	.m_data_3(\sdram|m_data[3]~q ),
	.m_data_4(\sdram|m_data[4]~q ),
	.m_data_5(\sdram|m_data[5]~q ),
	.m_data_6(\sdram|m_data[6]~q ),
	.m_data_7(\sdram|m_data[7]~q ),
	.m_data_8(\sdram|m_data[8]~q ),
	.m_data_9(\sdram|m_data[9]~q ),
	.m_data_10(\sdram|m_data[10]~q ),
	.m_data_11(\sdram|m_data[11]~q ),
	.m_data_12(\sdram|m_data[12]~q ),
	.m_data_13(\sdram|m_data[13]~q ),
	.m_data_14(\sdram|m_data[14]~q ),
	.m_data_15(\sdram|m_data[15]~q ),
	.m_data_16(\sdram|m_data[16]~q ),
	.m_data_17(\sdram|m_data[17]~q ),
	.m_data_18(\sdram|m_data[18]~q ),
	.m_data_19(\sdram|m_data[19]~q ),
	.m_data_20(\sdram|m_data[20]~q ),
	.m_data_21(\sdram|m_data[21]~q ),
	.m_data_22(\sdram|m_data[22]~q ),
	.m_data_23(\sdram|m_data[23]~q ),
	.m_data_24(\sdram|m_data[24]~q ),
	.m_data_25(\sdram|m_data[25]~q ),
	.m_data_26(\sdram|m_data[26]~q ),
	.m_data_27(\sdram|m_data[27]~q ),
	.m_data_28(\sdram|m_data[28]~q ),
	.m_data_29(\sdram|m_data[29]~q ),
	.m_data_30(\sdram|m_data[30]~q ),
	.m_data_31(\sdram|m_data[31]~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_22(\sdram|za_data[22]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_005|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_005|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_005|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_005|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_005|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_005|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_005|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_005|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_005|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_005|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_005|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_005|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_005|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_005|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_005|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_005|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_005|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_005|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_005|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_005|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_005|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_005|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_005|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_005|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_005|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_005|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_005|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_005|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_005|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_005|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_005|src_payload~31_combout ),
	.sdram_wire_dq_0(\sdram_wire_dq[0]~input_o ),
	.sdram_wire_dq_1(\sdram_wire_dq[1]~input_o ),
	.sdram_wire_dq_2(\sdram_wire_dq[2]~input_o ),
	.sdram_wire_dq_3(\sdram_wire_dq[3]~input_o ),
	.sdram_wire_dq_4(\sdram_wire_dq[4]~input_o ),
	.sdram_wire_dq_5(\sdram_wire_dq[5]~input_o ),
	.sdram_wire_dq_6(\sdram_wire_dq[6]~input_o ),
	.sdram_wire_dq_7(\sdram_wire_dq[7]~input_o ),
	.sdram_wire_dq_8(\sdram_wire_dq[8]~input_o ),
	.sdram_wire_dq_9(\sdram_wire_dq[9]~input_o ),
	.sdram_wire_dq_10(\sdram_wire_dq[10]~input_o ),
	.sdram_wire_dq_11(\sdram_wire_dq[11]~input_o ),
	.sdram_wire_dq_12(\sdram_wire_dq[12]~input_o ),
	.sdram_wire_dq_13(\sdram_wire_dq[13]~input_o ),
	.sdram_wire_dq_14(\sdram_wire_dq[14]~input_o ),
	.sdram_wire_dq_15(\sdram_wire_dq[15]~input_o ),
	.sdram_wire_dq_16(\sdram_wire_dq[16]~input_o ),
	.sdram_wire_dq_17(\sdram_wire_dq[17]~input_o ),
	.sdram_wire_dq_18(\sdram_wire_dq[18]~input_o ),
	.sdram_wire_dq_19(\sdram_wire_dq[19]~input_o ),
	.sdram_wire_dq_20(\sdram_wire_dq[20]~input_o ),
	.sdram_wire_dq_21(\sdram_wire_dq[21]~input_o ),
	.sdram_wire_dq_22(\sdram_wire_dq[22]~input_o ),
	.sdram_wire_dq_23(\sdram_wire_dq[23]~input_o ),
	.sdram_wire_dq_24(\sdram_wire_dq[24]~input_o ),
	.sdram_wire_dq_25(\sdram_wire_dq[25]~input_o ),
	.sdram_wire_dq_26(\sdram_wire_dq[26]~input_o ),
	.sdram_wire_dq_27(\sdram_wire_dq[27]~input_o ),
	.sdram_wire_dq_28(\sdram_wire_dq[28]~input_o ),
	.sdram_wire_dq_29(\sdram_wire_dq[29]~input_o ),
	.sdram_wire_dq_30(\sdram_wire_dq[30]~input_o ),
	.sdram_wire_dq_31(\sdram_wire_dq[31]~input_o ),
	.clk_clk(\clk_clk~input_o ));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .lut_mask = 64'hFFFBFFFFFFFEFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .shared_arith = "off";

assign \sdram_wire_dq[0]~input_o  = sdram_wire_dq[0];

assign \sdram_wire_dq[1]~input_o  = sdram_wire_dq[1];

assign \sdram_wire_dq[2]~input_o  = sdram_wire_dq[2];

assign \sdram_wire_dq[3]~input_o  = sdram_wire_dq[3];

assign \sdram_wire_dq[4]~input_o  = sdram_wire_dq[4];

assign \sdram_wire_dq[5]~input_o  = sdram_wire_dq[5];

assign \sdram_wire_dq[6]~input_o  = sdram_wire_dq[6];

assign \sdram_wire_dq[7]~input_o  = sdram_wire_dq[7];

assign \sdram_wire_dq[8]~input_o  = sdram_wire_dq[8];

assign \sdram_wire_dq[9]~input_o  = sdram_wire_dq[9];

assign \sdram_wire_dq[10]~input_o  = sdram_wire_dq[10];

assign \sdram_wire_dq[11]~input_o  = sdram_wire_dq[11];

assign \sdram_wire_dq[12]~input_o  = sdram_wire_dq[12];

assign \sdram_wire_dq[13]~input_o  = sdram_wire_dq[13];

assign \sdram_wire_dq[14]~input_o  = sdram_wire_dq[14];

assign \sdram_wire_dq[15]~input_o  = sdram_wire_dq[15];

assign \sdram_wire_dq[16]~input_o  = sdram_wire_dq[16];

assign \sdram_wire_dq[17]~input_o  = sdram_wire_dq[17];

assign \sdram_wire_dq[18]~input_o  = sdram_wire_dq[18];

assign \sdram_wire_dq[19]~input_o  = sdram_wire_dq[19];

assign \sdram_wire_dq[20]~input_o  = sdram_wire_dq[20];

assign \sdram_wire_dq[21]~input_o  = sdram_wire_dq[21];

assign \sdram_wire_dq[22]~input_o  = sdram_wire_dq[22];

assign \sdram_wire_dq[23]~input_o  = sdram_wire_dq[23];

assign \sdram_wire_dq[24]~input_o  = sdram_wire_dq[24];

assign \sdram_wire_dq[25]~input_o  = sdram_wire_dq[25];

assign \sdram_wire_dq[26]~input_o  = sdram_wire_dq[26];

assign \sdram_wire_dq[27]~input_o  = sdram_wire_dq[27];

assign \sdram_wire_dq[28]~input_o  = sdram_wire_dq[28];

assign \sdram_wire_dq[29]~input_o  = sdram_wire_dq[29];

assign \sdram_wire_dq[30]~input_o  = sdram_wire_dq[30];

assign \sdram_wire_dq[31]~input_o  = sdram_wire_dq[31];

assign \clk_clk~input_o  = clk_clk;

assign \sw_export[0]~input_o  = sw_export[0];

assign \sw_export[1]~input_o  = sw_export[1];

assign \sw_export[2]~input_o  = sw_export[2];

assign \sw_export[3]~input_o  = sw_export[3];

assign \sw_export[4]~input_o  = sw_export[4];

assign \sw_export[5]~input_o  = sw_export[5];

assign \sw_export[6]~input_o  = sw_export[6];

assign \sw_export[7]~input_o  = sw_export[7];

assign led_export[0] = \led|data_out[0]~q ;

assign led_export[1] = \led|data_out[1]~q ;

assign led_export[2] = \led|data_out[2]~q ;

assign led_export[3] = \led|data_out[3]~q ;

assign led_export[4] = \led|data_out[4]~q ;

assign led_export[5] = \led|data_out[5]~q ;

assign led_export[6] = \led|data_out[6]~q ;

assign led_export[7] = \led|data_out[7]~q ;

assign sdram_wire_addr[0] = \sdram|m_addr[0]~q ;

assign sdram_wire_addr[1] = \sdram|m_addr[1]~q ;

assign sdram_wire_addr[2] = \sdram|m_addr[2]~q ;

assign sdram_wire_addr[3] = \sdram|m_addr[3]~q ;

assign sdram_wire_addr[4] = \sdram|m_addr[4]~q ;

assign sdram_wire_addr[5] = \sdram|m_addr[5]~q ;

assign sdram_wire_addr[6] = \sdram|m_addr[6]~q ;

assign sdram_wire_addr[7] = \sdram|m_addr[7]~q ;

assign sdram_wire_addr[8] = \sdram|m_addr[8]~q ;

assign sdram_wire_addr[9] = \sdram|m_addr[9]~q ;

assign sdram_wire_addr[10] = \sdram|m_addr[10]~q ;

assign sdram_wire_addr[11] = \sdram|m_addr[11]~q ;

assign sdram_wire_addr[12] = \sdram|m_addr[12]~q ;

assign sdram_wire_ba[0] = \sdram|m_bank[0]~q ;

assign sdram_wire_ba[1] = \sdram|m_bank[1]~q ;

assign sdram_wire_cas_n = ~ \sdram|m_cmd[1]~q ;

assign sdram_wire_cke = vcc;

assign sdram_wire_cs_n = ~ \sdram|m_cmd[3]~q ;

assign sdram_wire_dqm[0] = \sdram|m_dqm[0]~q ;

assign sdram_wire_dqm[1] = \sdram|m_dqm[1]~q ;

assign sdram_wire_dqm[2] = \sdram|m_dqm[2]~q ;

assign sdram_wire_dqm[3] = \sdram|m_dqm[3]~q ;

assign sdram_wire_ras_n = ~ \sdram|m_cmd[2]~q ;

assign sdram_wire_we_n = ~ \sdram|m_cmd[0]~q ;

cyclonev_io_obuf \sdram_wire_dq[0]~output (
	.i(\sdram|m_data[0]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[0]),
	.obar());
defparam \sdram_wire_dq[0]~output .bus_hold = "false";
defparam \sdram_wire_dq[0]~output .open_drain_output = "false";
defparam \sdram_wire_dq[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[1]~output (
	.i(\sdram|m_data[1]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[1]),
	.obar());
defparam \sdram_wire_dq[1]~output .bus_hold = "false";
defparam \sdram_wire_dq[1]~output .open_drain_output = "false";
defparam \sdram_wire_dq[1]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[2]~output (
	.i(\sdram|m_data[2]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[2]),
	.obar());
defparam \sdram_wire_dq[2]~output .bus_hold = "false";
defparam \sdram_wire_dq[2]~output .open_drain_output = "false";
defparam \sdram_wire_dq[2]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[3]~output (
	.i(\sdram|m_data[3]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[3]),
	.obar());
defparam \sdram_wire_dq[3]~output .bus_hold = "false";
defparam \sdram_wire_dq[3]~output .open_drain_output = "false";
defparam \sdram_wire_dq[3]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[4]~output (
	.i(\sdram|m_data[4]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[4]),
	.obar());
defparam \sdram_wire_dq[4]~output .bus_hold = "false";
defparam \sdram_wire_dq[4]~output .open_drain_output = "false";
defparam \sdram_wire_dq[4]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[5]~output (
	.i(\sdram|m_data[5]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[5]),
	.obar());
defparam \sdram_wire_dq[5]~output .bus_hold = "false";
defparam \sdram_wire_dq[5]~output .open_drain_output = "false";
defparam \sdram_wire_dq[5]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[6]~output (
	.i(\sdram|m_data[6]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[6]),
	.obar());
defparam \sdram_wire_dq[6]~output .bus_hold = "false";
defparam \sdram_wire_dq[6]~output .open_drain_output = "false";
defparam \sdram_wire_dq[6]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[7]~output (
	.i(\sdram|m_data[7]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[7]),
	.obar());
defparam \sdram_wire_dq[7]~output .bus_hold = "false";
defparam \sdram_wire_dq[7]~output .open_drain_output = "false";
defparam \sdram_wire_dq[7]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[8]~output (
	.i(\sdram|m_data[8]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[8]),
	.obar());
defparam \sdram_wire_dq[8]~output .bus_hold = "false";
defparam \sdram_wire_dq[8]~output .open_drain_output = "false";
defparam \sdram_wire_dq[8]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[9]~output (
	.i(\sdram|m_data[9]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[9]),
	.obar());
defparam \sdram_wire_dq[9]~output .bus_hold = "false";
defparam \sdram_wire_dq[9]~output .open_drain_output = "false";
defparam \sdram_wire_dq[9]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[10]~output (
	.i(\sdram|m_data[10]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[10]),
	.obar());
defparam \sdram_wire_dq[10]~output .bus_hold = "false";
defparam \sdram_wire_dq[10]~output .open_drain_output = "false";
defparam \sdram_wire_dq[10]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[11]~output (
	.i(\sdram|m_data[11]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[11]),
	.obar());
defparam \sdram_wire_dq[11]~output .bus_hold = "false";
defparam \sdram_wire_dq[11]~output .open_drain_output = "false";
defparam \sdram_wire_dq[11]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[12]~output (
	.i(\sdram|m_data[12]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[12]),
	.obar());
defparam \sdram_wire_dq[12]~output .bus_hold = "false";
defparam \sdram_wire_dq[12]~output .open_drain_output = "false";
defparam \sdram_wire_dq[12]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[13]~output (
	.i(\sdram|m_data[13]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[13]),
	.obar());
defparam \sdram_wire_dq[13]~output .bus_hold = "false";
defparam \sdram_wire_dq[13]~output .open_drain_output = "false";
defparam \sdram_wire_dq[13]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[14]~output (
	.i(\sdram|m_data[14]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[14]),
	.obar());
defparam \sdram_wire_dq[14]~output .bus_hold = "false";
defparam \sdram_wire_dq[14]~output .open_drain_output = "false";
defparam \sdram_wire_dq[14]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[15]~output (
	.i(\sdram|m_data[15]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[15]),
	.obar());
defparam \sdram_wire_dq[15]~output .bus_hold = "false";
defparam \sdram_wire_dq[15]~output .open_drain_output = "false";
defparam \sdram_wire_dq[15]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[16]~output (
	.i(\sdram|m_data[16]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[16]),
	.obar());
defparam \sdram_wire_dq[16]~output .bus_hold = "false";
defparam \sdram_wire_dq[16]~output .open_drain_output = "false";
defparam \sdram_wire_dq[16]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[17]~output (
	.i(\sdram|m_data[17]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[17]),
	.obar());
defparam \sdram_wire_dq[17]~output .bus_hold = "false";
defparam \sdram_wire_dq[17]~output .open_drain_output = "false";
defparam \sdram_wire_dq[17]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[18]~output (
	.i(\sdram|m_data[18]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[18]),
	.obar());
defparam \sdram_wire_dq[18]~output .bus_hold = "false";
defparam \sdram_wire_dq[18]~output .open_drain_output = "false";
defparam \sdram_wire_dq[18]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[19]~output (
	.i(\sdram|m_data[19]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[19]),
	.obar());
defparam \sdram_wire_dq[19]~output .bus_hold = "false";
defparam \sdram_wire_dq[19]~output .open_drain_output = "false";
defparam \sdram_wire_dq[19]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[20]~output (
	.i(\sdram|m_data[20]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[20]),
	.obar());
defparam \sdram_wire_dq[20]~output .bus_hold = "false";
defparam \sdram_wire_dq[20]~output .open_drain_output = "false";
defparam \sdram_wire_dq[20]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[21]~output (
	.i(\sdram|m_data[21]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[21]),
	.obar());
defparam \sdram_wire_dq[21]~output .bus_hold = "false";
defparam \sdram_wire_dq[21]~output .open_drain_output = "false";
defparam \sdram_wire_dq[21]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[22]~output (
	.i(\sdram|m_data[22]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[22]),
	.obar());
defparam \sdram_wire_dq[22]~output .bus_hold = "false";
defparam \sdram_wire_dq[22]~output .open_drain_output = "false";
defparam \sdram_wire_dq[22]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[23]~output (
	.i(\sdram|m_data[23]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[23]),
	.obar());
defparam \sdram_wire_dq[23]~output .bus_hold = "false";
defparam \sdram_wire_dq[23]~output .open_drain_output = "false";
defparam \sdram_wire_dq[23]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[24]~output (
	.i(\sdram|m_data[24]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[24]),
	.obar());
defparam \sdram_wire_dq[24]~output .bus_hold = "false";
defparam \sdram_wire_dq[24]~output .open_drain_output = "false";
defparam \sdram_wire_dq[24]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[25]~output (
	.i(\sdram|m_data[25]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[25]),
	.obar());
defparam \sdram_wire_dq[25]~output .bus_hold = "false";
defparam \sdram_wire_dq[25]~output .open_drain_output = "false";
defparam \sdram_wire_dq[25]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[26]~output (
	.i(\sdram|m_data[26]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[26]),
	.obar());
defparam \sdram_wire_dq[26]~output .bus_hold = "false";
defparam \sdram_wire_dq[26]~output .open_drain_output = "false";
defparam \sdram_wire_dq[26]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[27]~output (
	.i(\sdram|m_data[27]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[27]),
	.obar());
defparam \sdram_wire_dq[27]~output .bus_hold = "false";
defparam \sdram_wire_dq[27]~output .open_drain_output = "false";
defparam \sdram_wire_dq[27]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[28]~output (
	.i(\sdram|m_data[28]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[28]),
	.obar());
defparam \sdram_wire_dq[28]~output .bus_hold = "false";
defparam \sdram_wire_dq[28]~output .open_drain_output = "false";
defparam \sdram_wire_dq[28]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[29]~output (
	.i(\sdram|m_data[29]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[29]),
	.obar());
defparam \sdram_wire_dq[29]~output .bus_hold = "false";
defparam \sdram_wire_dq[29]~output .open_drain_output = "false";
defparam \sdram_wire_dq[29]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[30]~output (
	.i(\sdram|m_data[30]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[30]),
	.obar());
defparam \sdram_wire_dq[30]~output .bus_hold = "false";
defparam \sdram_wire_dq[30]~output .open_drain_output = "false";
defparam \sdram_wire_dq[30]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \sdram_wire_dq[31]~output (
	.i(\sdram|m_data[31]~q ),
	.oe(\sdram|oe~q ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[31]),
	.obar());
defparam \sdram_wire_dq[31]~output .bus_hold = "false";
defparam \sdram_wire_dq[31]~output .open_drain_output = "false";
defparam \sdram_wire_dq[31]~output .shift_series_termination_control = "false";

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .lut_mask = 64'hF3FFFFFF77FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 64'hFDF7FFFFF7FDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'hF9FFF6FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hFF7FFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|ir_out[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h7DD77DD7D77DD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\nios2|cpu|the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_tck|sr[0]~q ),
	.datad(!\jtag_uart|sdram_demo_jtag_uart_alt_jtag_atlantic|adapted_tdo~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFAAAAFFAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hFBFEFEFBFEFBFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hAAFFFFAAAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFFFDF8FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hBFFFBF3FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module sdram_demo_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	resetrequest,
	altera_reset_synchronizer_int_chain_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
input 	resetrequest;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


sdram_demo_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

sdram_demo_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.resetrequest(resetrequest),
	.clk(clk_clk));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module sdram_demo_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	resetrequest,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	resetrequest;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module sdram_demo_sdram_demo_jtag_uart (
	W_alu_result_2,
	d_writedata_10,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	adapted_tdo,
	d_writedata_0,
	r_sync_rst,
	always0,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	av_begintransfer,
	Equal5,
	av_waitrequest1,
	mem_used_1,
	read_latency_shift_reg,
	b_full,
	ien_AF1,
	read_01,
	ien_AE1,
	av_readdata_9,
	av_readdata_8,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	b_full1,
	rvalid1,
	woverflow1,
	ac1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	d_writedata_10;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	Add1;
output 	Add11;
output 	Add12;
output 	Add13;
output 	Add14;
output 	Add15;
output 	Add16;
output 	adapted_tdo;
input 	d_writedata_0;
input 	r_sync_rst;
input 	always0;
output 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	av_begintransfer;
input 	Equal5;
output 	av_waitrequest1;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full;
output 	ien_AF1;
output 	read_01;
output 	ien_AE1;
output 	av_readdata_9;
output 	av_readdata_8;
output 	b_non_empty;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	b_full1;
output 	rvalid1;
output 	woverflow1;
output 	ac1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|r_ena1~q ;
wire \fifo_wr~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \rvalid~0_combout ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|t_ena~reg0_q ;
wire \wr_rfifo~combout ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[0]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|t_pause~reg0_q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[1]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[2]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[3]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[4]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[5]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[6]~q ;
wire \sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[7]~q ;
wire \fifo_wr~0_combout ;
wire \Add1~2 ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \Add1~26 ;
wire \av_waitrequest~0_combout ;
wire \ien_AE~0_combout ;
wire \fifo_rd~0_combout ;
wire \fifo_rd~1_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \fifo_AF~q ;
wire \rvalid~1_combout ;
wire \woverflow~0_combout ;
wire \ac~0_combout ;


sdram_demo_sdram_demo_jtag_uart_scfifo_w the_sdram_demo_jtag_uart_scfifo_w(
	.q_b_7(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.fifo_wr(\fifo_wr~q ),
	.b_non_empty(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.b_full(b_full1),
	.counter_reg_bit_3(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_5(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_jtag_uart_scfifo_r the_sdram_demo_jtag_uart_scfifo_r(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.r_sync_rst(r_sync_rst),
	.Equal5(Equal5),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(\fifo_rd~0_combout ),
	.rvalid(\rvalid~0_combout ),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(\sdram_demo_jtag_uart_alt_jtag_atlantic|t_ena~reg0_q ),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

sdram_demo_alt_jtag_atlantic sdram_demo_jtag_uart_alt_jtag_atlantic(
	.r_dat({\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.adapted_tdo1(adapted_tdo),
	.rst_n(r_sync_rst),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\sdram_demo_jtag_uart_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\sdram_demo_jtag_uart_alt_jtag_atlantic|r_ena1~q ),
	.t_ena(\sdram_demo_jtag_uart_alt_jtag_atlantic|t_ena~reg0_q ),
	.wdata_0(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.t_pause(\sdram_demo_jtag_uart_alt_jtag_atlantic|t_pause~reg0_q ),
	.wdata_1(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\sdram_demo_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \r_val~0 (
	.dataa(!\sdram_demo_jtag_uart_alt_jtag_atlantic|rvalid0~q ),
	.datab(!\r_val~q ),
	.datac(!\sdram_demo_jtag_uart_alt_jtag_atlantic|r_ena1~q ),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_val~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_val~0 .extended_lut = "off";
defparam \r_val~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \r_val~0 .shared_arith = "off";

cyclonev_lcell_comb \rvalid~0 (
	.dataa(!Equal5),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg),
	.datad(!b_non_empty),
	.datae(!\fifo_rd~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~0 .extended_lut = "off";
defparam \rvalid~0 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \rvalid~0 .shared_arith = "off";

cyclonev_lcell_comb wr_rfifo(
	.dataa(!b_full),
	.datab(!\sdram_demo_jtag_uart_alt_jtag_atlantic|t_ena~reg0_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_rfifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wr_rfifo.extended_lut = "off";
defparam wr_rfifo.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam wr_rfifo.shared_arith = "off";

cyclonev_lcell_comb \fifo_wr~0 (
	.dataa(!W_alu_result_2),
	.datab(!always0),
	.datac(!\av_waitrequest~0_combout ),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr~0 .extended_lut = "off";
defparam \fifo_wr~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \fifo_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add1),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add11),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add12),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add13),
	.cout(),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add14),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add15),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add16),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AF1),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AE1),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclonev_lcell_comb \av_readdata[9] (
	.dataa(!\fifo_AE~q ),
	.datab(!ien_AE1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[9] .extended_lut = "off";
defparam \av_readdata[9] .lut_mask = 64'h7777777777777777;
defparam \av_readdata[9] .shared_arith = "off";

cyclonev_lcell_comb \av_readdata[8]~0 (
	.dataa(!ien_AF1),
	.datab(!\pause_irq~q ),
	.datac(!\fifo_AF~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[8]~0 .extended_lut = "off";
defparam \av_readdata[8]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_readdata[8]~0 .shared_arith = "off";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!av_begintransfer),
	.datab(!Equal5),
	.datac(!av_waitrequest1),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \av_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \ien_AE~0 (
	.dataa(!W_alu_result_2),
	.datab(!always0),
	.datac(!av_begintransfer),
	.datad(!Equal5),
	.datae(!av_waitrequest1),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ien_AE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ien_AE~0 .extended_lut = "off";
defparam \ien_AE~0 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \ien_AE~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~0 (
	.dataa(!W_alu_result_2),
	.datab(!av_waitrequest1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~0 .extended_lut = "off";
defparam \fifo_rd~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \fifo_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~1 (
	.dataa(!Equal5),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg),
	.datad(!\fifo_rd~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~1 .extended_lut = "off";
defparam \fifo_rd~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \fifo_rd~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datab(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datac(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!b_full1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datad(!\the_sdram_demo_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cyclonev_lcell_comb \pause_irq~0 (
	.dataa(!read_01),
	.datab(!\pause_irq~q ),
	.datac(!b_non_empty),
	.datad(!\sdram_demo_jtag_uart_alt_jtag_atlantic|t_pause~reg0_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pause_irq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pause_irq~0 .extended_lut = "off";
defparam \pause_irq~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \pause_irq~0 .shared_arith = "off";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(!counter_reg_bit_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000000000000000;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add0~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add0~9_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan1~1 .shared_arith = "off";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclonev_lcell_comb \rvalid~1 (
	.dataa(!b_non_empty),
	.datab(!\fifo_rd~1_combout ),
	.datac(!rvalid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~1 .extended_lut = "off";
defparam \rvalid~1 .lut_mask = 64'h4747474747474747;
defparam \rvalid~1 .shared_arith = "off";

cyclonev_lcell_comb \woverflow~0 (
	.dataa(!W_alu_result_2),
	.datab(!always0),
	.datac(!\av_waitrequest~0_combout ),
	.datad(!b_full1),
	.datae(!woverflow1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~0 .extended_lut = "off";
defparam \woverflow~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \woverflow~0 .shared_arith = "off";

cyclonev_lcell_comb \ac~0 (
	.dataa(!d_writedata_10),
	.datab(!\sdram_demo_jtag_uart_alt_jtag_atlantic|t_ena~reg0_q ),
	.datac(!\ien_AE~0_combout ),
	.datad(!\sdram_demo_jtag_uart_alt_jtag_atlantic|t_pause~reg0_q ),
	.datae(!ac1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac~0 .extended_lut = "off";
defparam \ac~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ac~0 .shared_arith = "off";

endmodule

module sdram_demo_alt_jtag_atlantic (
	r_dat,
	adapted_tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_ena,
	wdata_0,
	t_pause,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	adapted_tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_ena;
output 	wdata_0;
output 	t_pause;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state~1_combout ;
wire \state~q ;
wire \td_shift[0]~2_combout ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[4]~q ;
wire \count[5]~q ;
wire \count[6]~q ;
wire \count[7]~q ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count[9]~_wirecell_combout ;
wire \count[0]~q ;
wire \count[1]~q ;
wire \state~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~3_combout ;
wire \td_shift[9]~q ;
wire \td_shift~0_combout ;
wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~q ;
wire \td_shift~4_combout ;
wire \rdata[0]~q ;
wire \rdata[6]~q ;
wire \td_shift~12_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~11_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~10_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~9_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~8_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~7_combout ;
wire \td_shift[3]~q ;
wire \td_shift~6_combout ;
wire \td_shift[2]~q ;
wire \td_shift~5_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~1_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read_req~q ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \rst2~q ;
wire \rvalid0~1_combout ;
wire \write~0_combout ;
wire \wdata[1]~0_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~0_combout ;
wire \write_valid~q ;
wire \t_ena~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \always2~1_combout ;
wire \t_pause~0_combout ;


dffeas adapted_tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(adapted_tdo1),
	.prn(vcc));
defparam adapted_tdo.is_wysiwyg = "true";
defparam adapted_tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas \t_ena~reg0 (
	.clk(clk),
	.d(\t_ena~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena),
	.prn(vcc));
defparam \t_ena~reg0 .is_wysiwyg = "true";
defparam \t_ena~reg0 .power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \t_pause~reg0 (
	.clk(clk),
	.d(\t_pause~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause),
	.prn(vcc));
defparam \t_pause~reg0 .is_wysiwyg = "true";
defparam \t_pause~reg0 .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cyclonev_lcell_comb \state~1 (
	.dataa(!splitter_nodes_receive_0_3),
	.datab(!virtual_ir_scan_reg),
	.datac(!state_3),
	.datad(!state_4),
	.datae(!\state~q ),
	.dataf(!altera_internal_jtag1),
	.datag(!irf_reg_0_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~1 .extended_lut = "on";
defparam \state~1 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \state~1 .shared_arith = "off";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclonev_lcell_comb \td_shift[0]~2 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift[0]~2 .extended_lut = "off";
defparam \td_shift[0]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \td_shift[0]~2 .shared_arith = "off";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclonev_lcell_comb \count[9]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!altera_internal_jtag1),
	.datad(!state_4),
	.datae(!\count[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~0 .extended_lut = "off";
defparam \count[9]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \count[9]~0 .shared_arith = "off";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclonev_lcell_comb \count[9]~_wirecell (
	.dataa(!\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~_wirecell .extended_lut = "off";
defparam \count[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count[9]~_wirecell .shared_arith = "off";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count[9]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \state~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \state~0 .shared_arith = "off";

cyclonev_lcell_comb \user_saw_rvalid~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\td_shift[0]~q ),
	.datac(!\state~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\state~0_combout ),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_saw_rvalid~0 .extended_lut = "off";
defparam \user_saw_rvalid~0 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \user_saw_rvalid~0 .shared_arith = "off";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cyclonev_lcell_comb \r_ena~0 (
	.dataa(!r_val),
	.datab(!r_ena11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_ena~0 .extended_lut = "off";
defparam \r_ena~0 .lut_mask = 64'h7777777777777777;
defparam \r_ena~0 .shared_arith = "off";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~3 (
	.dataa(!\count[9]~q ),
	.datab(!\td_shift[10]~q ),
	.datac(!\rdata[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~3 .extended_lut = "off";
defparam \td_shift~3 .lut_mask = 64'h2727272727272727;
defparam \td_shift~3 .shared_arith = "off";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclonev_lcell_comb \td_shift~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~0 .extended_lut = "off";
defparam \td_shift~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \td_shift~0 .shared_arith = "off";

cyclonev_lcell_comb \tck_t_dav~0 (
	.dataa(!t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tck_t_dav~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tck_t_dav~0 .extended_lut = "off";
defparam \tck_t_dav~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \tck_t_dav~0 .shared_arith = "off";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclonev_lcell_comb \write_stalled~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\tck_t_dav~q ),
	.datac(!\td_shift[10]~q ),
	.datad(!\write_stalled~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~0 .extended_lut = "off";
defparam \write_stalled~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \write_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \write_stalled~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!state_4),
	.datae(!virtual_ir_scan_reg),
	.dataf(!splitter_nodes_receive_0_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~1 .extended_lut = "off";
defparam \write_stalled~1 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \write_stalled~1 .shared_arith = "off";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclonev_lcell_comb \td_shift~4 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~4 .extended_lut = "off";
defparam \td_shift~4 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \td_shift~4 .shared_arith = "off";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~12 (
	.dataa(!\td_shift[9]~q ),
	.datab(!\count[9]~q ),
	.datac(!\rdata[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~12 .extended_lut = "off";
defparam \td_shift~12 .lut_mask = 64'h4747474747474747;
defparam \td_shift~12 .shared_arith = "off";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclonev_lcell_comb \td_shift~11 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[8]~q ),
	.datae(!\rdata[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~11 .extended_lut = "off";
defparam \td_shift~11 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~11 .shared_arith = "off";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cyclonev_lcell_comb \td_shift~10 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[7]~q ),
	.dataf(!\rdata[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~10 .extended_lut = "off";
defparam \td_shift~10 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~10 .shared_arith = "off";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~9 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[6]~q ),
	.dataf(!\rdata[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~9 .extended_lut = "off";
defparam \td_shift~9 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~9 .shared_arith = "off";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~8 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[5]~q ),
	.datae(!\rdata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~8 .extended_lut = "off";
defparam \td_shift~8 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~8 .shared_arith = "off";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclonev_lcell_comb \td_shift~7 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[4]~q ),
	.datae(!\rdata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~7 .extended_lut = "off";
defparam \td_shift~7 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~7 .shared_arith = "off";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~6 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[0]~q ),
	.dataf(!\td_shift[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~6 .extended_lut = "off";
defparam \td_shift~6 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~6 .shared_arith = "off";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~5 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\write_stalled~q ),
	.datae(!\td_shift~4_combout ),
	.dataf(!\td_shift[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~5 .extended_lut = "off";
defparam \td_shift~5 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \td_shift~5 .shared_arith = "off";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \td_shift~1 (
	.dataa(!\state~q ),
	.datab(!\td_shift~0_combout ),
	.datac(!\tck_t_dav~q ),
	.datad(!\td_shift[1]~q ),
	.datae(!\count[9]~q ),
	.dataf(!\rvalid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~1 .extended_lut = "off";
defparam \td_shift~1 .lut_mask = 64'hBFFFEFFFFFFFFFFF;
defparam \td_shift~1 .shared_arith = "off";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclonev_lcell_comb \rvalid0~0 (
	.dataa(!rvalid01),
	.datab(!r_val),
	.datac(!r_ena11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~0 .extended_lut = "off";
defparam \rvalid0~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \rvalid0~0 .shared_arith = "off";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \read~0 .shared_arith = "off";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclonev_lcell_comb \rvalid0~1 (
	.dataa(!\user_saw_rvalid~q ),
	.datab(!\rvalid0~0_combout ),
	.datac(!\read_req~q ),
	.datad(!\read1~q ),
	.datae(!\read2~q ),
	.dataf(!\rst2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~1 .extended_lut = "off";
defparam \rvalid0~1 .lut_mask = 64'hFFFFFFFFFEFFFFFE;
defparam \rvalid0~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \wdata[1]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!state_4),
	.datad(!virtual_ir_scan_reg),
	.datae(!splitter_nodes_receive_0_3),
	.dataf(!\count[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata[1]~0 .extended_lut = "off";
defparam \wdata[1]~0 .lut_mask = 64'hFFBFFFFFFFFFFFFF;
defparam \wdata[1]~0 .shared_arith = "off";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\write1~q ),
	.datab(!\write2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h6666666666666666;
defparam \always2~0 .shared_arith = "off";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclonev_lcell_comb \t_ena~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!t_ena),
	.datae(!\always2~0_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_ena~0 .extended_lut = "off";
defparam \t_ena~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \t_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \jupdate~0 (
	.dataa(!irf_reg_0_1),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!\jupdate~q ),
	.datae(!state_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jupdate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jupdate~0 .extended_lut = "off";
defparam \jupdate~0 .lut_mask = 64'h9669699696696996;
defparam \jupdate~0 .shared_arith = "off";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\jupdate1~q ),
	.datab(!\jupdate2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h6666666666666666;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \t_pause~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!\always2~0_combout ),
	.datae(!\write_valid~q ),
	.dataf(!\always2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_pause~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_pause~0 .extended_lut = "off";
defparam \t_pause~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \t_pause~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_jtag_uart_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	Equal5,
	mem_used_1,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	rvalid,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
input 	Equal5;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	rvalid;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.Equal5(Equal5),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.rvalid(rvalid),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module sdram_demo_scfifo_1 (
	q,
	r_sync_rst,
	Equal5,
	mem_used_1,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	rvalid,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	Equal5;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	rvalid;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_scfifo_3291 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.Equal5(Equal5),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.rvalid(rvalid),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module sdram_demo_scfifo_3291 (
	q,
	r_sync_rst,
	Equal5,
	mem_used_1,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	rvalid,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	Equal5;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	rvalid;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_a_dpfifo_5771 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.Equal5(Equal5),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.rvalid(rvalid),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module sdram_demo_a_dpfifo_5771 (
	q,
	r_sync_rst,
	Equal5,
	mem_used_1,
	read_latency_shift_reg,
	b_full,
	b_non_empty,
	fifo_rd,
	rvalid,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	Equal5;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	rvalid;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


sdram_demo_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.Equal5(Equal5),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.fifo_rd(fifo_rd),
	.rvalid(rvalid),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wreq),
	.clock(clock));

sdram_demo_cntr_jgb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

sdram_demo_cntr_jgb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.rvalid(rvalid),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

sdram_demo_altsyncram_7pu1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(rvalid),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

endmodule

module sdram_demo_a_fefifo_7cf (
	r_sync_rst,
	Equal5,
	mem_used_1,
	read_latency_shift_reg,
	b_full1,
	b_non_empty1,
	fifo_rd,
	rvalid,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	Equal5;
input 	mem_used_1;
input 	read_latency_shift_reg;
output 	b_full1;
output 	b_non_empty1;
input 	fifo_rd;
input 	rvalid;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \b_non_empty~0_combout ;


sdram_demo_cntr_vg7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wr_rfifo),
	._(\_~2_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~2 (
	.dataa(!Equal5),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg),
	.datad(!b_non_empty1),
	.datae(!fifo_rd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h6996966996696996;
defparam \_~2 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!b_non_empty1),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!counter_reg_bit_3),
	.datae(!counter_reg_bit_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!rvalid),
	.datac(!counter_reg_bit_1),
	.datad(!counter_reg_bit_0),
	.datae(!t_ena),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \_~0 (
	.dataa(!counter_reg_bit_5),
	.datab(!counter_reg_bit_4),
	.datac(!counter_reg_bit_3),
	.datad(!wr_rfifo),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \_~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_0),
	.datad(!\_~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!b_full1),
	.datab(!b_non_empty1),
	.datac(!rvalid),
	.datad(!t_ena),
	.datae(!\_~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hF7FFD5FFF7FFD5FF;
defparam \b_non_empty~0 .shared_arith = "off";

endmodule

module sdram_demo_cntr_vg7 (
	r_sync_rst,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_altsyncram_7pu1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_r:the_sdram_demo_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module sdram_demo_cntr_jgb (
	r_sync_rst,
	rvalid,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	rvalid;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_cntr_jgb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_jtag_uart_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	fifo_wr,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	fifo_wr;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.wrreq(fifo_wr),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clk_clk));

endmodule

module sdram_demo_scfifo_2 (
	q,
	data,
	r_sync_rst,
	wrreq,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wrreq;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_scfifo_3291_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.wrreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module sdram_demo_scfifo_3291_1 (
	q,
	data,
	r_sync_rst,
	wrreq,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wrreq;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_a_dpfifo_5771_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.wreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.b_full(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module sdram_demo_a_dpfifo_5771_1 (
	q,
	data,
	r_sync_rst,
	wreq,
	b_non_empty,
	r_val,
	b_full,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	wreq;
output 	b_non_empty;
input 	r_val;
output 	b_full;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


sdram_demo_altsyncram_7pu1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.clocken1(r_val),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

sdram_demo_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.b_full1(b_full),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

sdram_demo_cntr_jgb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

sdram_demo_cntr_jgb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

endmodule

module sdram_demo_a_fefifo_7cf_1 (
	r_sync_rst,
	fifo_wr,
	b_non_empty1,
	r_val,
	b_full1,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	b_non_empty1;
input 	r_val;
output 	b_full1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;


sdram_demo_cntr_vg7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(fifo_wr),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!fifo_wr),
	.datab(!r_val),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h6666666666666666;
defparam \_~0 .shared_arith = "off";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \b_non_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~1 (
	.dataa(!r_val),
	.datab(!counter_reg_bit_3),
	.datac(!counter_reg_bit_0),
	.datad(!\b_non_empty~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~1 .extended_lut = "off";
defparam \b_non_empty~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \b_non_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~2 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!b_full1),
	.datad(!\b_non_empty~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~2 .extended_lut = "off";
defparam \b_non_empty~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \b_non_empty~2 .shared_arith = "off";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_5),
	.datae(!counter_reg_bit_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!r_val),
	.datab(!b_full1),
	.datac(!counter_reg_bit_0),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_1),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

endmodule

module sdram_demo_cntr_vg7_1 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_altsyncram_7pu1_1 (
	q_b,
	data_a,
	wren_a,
	clocken1,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	wren_a;
input 	clocken1;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "sdram_demo_jtag_uart:jtag_uart|sdram_demo_jtag_uart_scfifo_w:the_sdram_demo_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module sdram_demo_cntr_jgb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_cntr_jgb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_led (
	W_alu_result_4,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	reset_n,
	d_write,
	write_accepted,
	always0,
	Equal4,
	rst1,
	wait_latency_counter_1,
	always01,
	wait_latency_counter_0,
	mem_used_1,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	reset_n;
input 	d_write;
input 	write_accepted;
output 	always0;
input 	Equal4;
input 	rst1;
input 	wait_latency_counter_1;
output 	always01;
input 	wait_latency_counter_0;
input 	mem_used_1;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~2_combout ;
wire \always0~3_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!d_write),
	.datab(!write_accepted),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always0),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!rst1),
	.datab(!wait_latency_counter_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always01),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!W_alu_result_2),
	.datac(!W_alu_result_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \always0~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!mem_used_1),
	.datac(!W_alu_result_2),
	.datad(!W_alu_result_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~2 .extended_lut = "off";
defparam \always0~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \always0~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~3 (
	.dataa(!always0),
	.datab(!W_alu_result_4),
	.datac(!Equal4),
	.datad(!always01),
	.datae(!\always0~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~3 .extended_lut = "off";
defparam \always0~3 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always0~3 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_24,
	W_alu_result_25,
	W_alu_result_26,
	W_alu_result_27,
	W_alu_result_28,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_21,
	W_alu_result_22,
	W_alu_result_23,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_17,
	F_pc_16,
	F_pc_18,
	F_pc_19,
	F_pc_20,
	F_pc_21,
	F_pc_22,
	F_pc_23,
	F_pc_24,
	F_pc_26,
	F_pc_15,
	F_pc_14,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	ram_block1a32,
	ram_block1a0,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a37,
	ram_block1a5,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	readdata_0,
	q_b_0,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_5,
	readdata_8,
	readdata_10,
	readdata_9,
	readdata_28,
	readdata_21,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_17,
	readdata_18,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_21,
	av_readdata_pre_22,
	readdata_27,
	av_readdata_pre_18,
	av_readdata_pre_17,
	readdata_7,
	readdata_6,
	av_readdata_pre_16,
	readdata_20,
	readdata_19,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	d_writedata_0,
	r_sync_rst,
	d_write,
	write_accepted,
	always0,
	Equal4,
	rst1,
	wait_latency_counter_1,
	always01,
	wait_latency_counter_0,
	mem_used_1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	entries_1,
	entries_0,
	d_read,
	nios2_data_master_waitrequest,
	av_begintransfer,
	sink_ready,
	saved_grant_0,
	WideOr0,
	saved_grant_01,
	mem_used_11,
	Equal5,
	saved_grant_02,
	waitrequest,
	mem_used_12,
	av_waitrequest,
	mem_used_13,
	WideOr01,
	src0_valid,
	za_valid,
	src0_valid1,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	av_waitrequest1,
	Equal1,
	src5_valid,
	saved_grant_1,
	i_read,
	F_pc_25,
	src_valid,
	src_data_68,
	src_data_58,
	src_valid1,
	src_data_59,
	src_data_60,
	src_data_61,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_50,
	src_data_51,
	m0_write,
	m0_write1,
	src_data_52,
	src_data_53,
	src_data_54,
	src_data_55,
	src_data_56,
	src_data_57,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	src_valid2,
	rf_source_valid,
	read_latency_shift_reg,
	src1_valid,
	src1_valid1,
	src1_valid2,
	WideOr12,
	hbreak_enabled,
	src0_valid2,
	av_readdata_pre_0,
	za_data_0,
	address_reg_a_0,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	za_data_24,
	av_readdata_pre_24,
	za_data_25,
	av_readdata_pre_25,
	za_data_26,
	av_readdata_pre_26,
	za_data_1,
	av_readdata_pre_1,
	za_data_4,
	av_readdata_pre_4,
	za_data_3,
	av_readdata_pre_3,
	za_data_2,
	av_readdata_pre_2,
	WideOr13,
	src_data_461,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_161,
	za_data_5,
	av_readdata_pre_5,
	av_readdata_pre_8,
	av_readdata_pre_10,
	av_readdata_pre_9,
	za_data_28,
	av_readdata_pre_28,
	av_readdata_pre_211,
	za_data_29,
	av_readdata_pre_29,
	za_data_30,
	av_readdata_pre_30,
	za_data_31,
	av_readdata_pre_31,
	av_readdata_pre_171,
	av_readdata_pre_181,
	za_data_27,
	av_readdata_pre_27,
	za_data_7,
	av_readdata_pre_7,
	za_data_6,
	av_readdata_pre_6,
	av_readdata_pre_201,
	av_readdata_pre_191,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	b_full,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	d_writedata_24,
	src_payload24,
	d_writedata_25,
	src_payload25,
	d_writedata_26,
	src_payload26,
	d_writedata_27,
	src_payload27,
	d_writedata_28,
	src_payload28,
	d_writedata_29,
	src_payload29,
	d_writedata_30,
	src_payload30,
	d_writedata_31,
	src_payload31,
	readdata_01,
	src_data_511,
	src_payload32,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_462,
	src_data_471,
	src_data_481,
	src_data_491,
	src_data_501,
	src_data_32,
	ien_AF,
	read_0,
	readdata_02,
	av_readdata_pre_81,
	ien_AE,
	av_readdata_9,
	av_readdata_8,
	src_payload33,
	src_data_34,
	src_payload34,
	src_payload35,
	src_data_35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_data_33,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	src_payload51,
	av_readdata_pre_91,
	src_payload52,
	src_data_24,
	src_payload53,
	src_payload54,
	src_data_25,
	src_payload55,
	src_data_26,
	src_payload56,
	src_data_27,
	src_payload57,
	src_data_28,
	src_payload58,
	src_payload59,
	src_payload60,
	src_payload61,
	src_payload62,
	av_readdata_pre_151,
	src_payload63,
	av_readdata_pre_141,
	av_readdata_pre_131,
	av_readdata_pre_121,
	av_readdata_pre_101,
	readdata_110,
	readdata_111,
	readdata_210,
	readdata_211,
	readdata_32,
	readdata_33,
	readdata_41,
	readdata_42,
	readdata_51,
	readdata_52,
	readdata_61,
	readdata_62,
	readdata_71,
	readdata_72,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	src_payload64,
	src_data_382,
	src_data_402,
	src_data_392,
	src_data_452,
	src_data_442,
	src_data_432,
	src_data_422,
	src_data_412,
	src_payload65,
	src_data_321,
	b_full1,
	src_data_29,
	src_data_30,
	src_data_31,
	rvalid,
	woverflow,
	ac,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_data_341,
	src_payload70,
	src_payload71,
	src_data_351,
	src_payload72,
	src_payload73,
	src_payload74,
	src_payload75,
	src_data_331,
	src_payload76,
	src_payload77,
	src_payload78,
	src_payload79,
	src_payload80,
	src_payload81,
	src_payload82,
	src_payload83,
	src_payload84,
	src_payload85,
	src_payload86,
	src_payload87,
	src_payload88,
	src_payload89,
	src_payload90,
	src_payload91,
	src_payload92,
	src_payload93,
	src_payload94,
	src_payload95,
	src_payload96,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_9;
input 	W_alu_result_24;
input 	W_alu_result_25;
input 	W_alu_result_26;
input 	W_alu_result_27;
input 	W_alu_result_28;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_21;
input 	W_alu_result_22;
input 	W_alu_result_23;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_8;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_18;
input 	F_pc_19;
input 	F_pc_20;
input 	F_pc_21;
input 	F_pc_22;
input 	F_pc_23;
input 	F_pc_24;
input 	F_pc_26;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_9;
input 	F_pc_11;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_10;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
input 	F_pc_8;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a38;
input 	ram_block1a6;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	readdata_0;
input 	q_b_0;
input 	readdata_22;
input 	readdata_23;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_1;
input 	readdata_4;
input 	readdata_3;
input 	readdata_2;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	readdata_14;
input 	readdata_15;
input 	readdata_16;
input 	readdata_5;
input 	readdata_8;
input 	readdata_10;
input 	readdata_9;
input 	readdata_28;
input 	readdata_21;
input 	readdata_29;
input 	readdata_30;
input 	readdata_31;
input 	readdata_17;
input 	readdata_18;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
input 	readdata_27;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
input 	readdata_7;
input 	readdata_6;
output 	av_readdata_pre_16;
input 	readdata_20;
input 	readdata_19;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	Add1;
input 	Add11;
input 	Add12;
input 	Add13;
input 	Add14;
input 	Add15;
input 	Add16;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_write;
output 	write_accepted;
input 	always0;
output 	Equal4;
input 	rst1;
output 	wait_latency_counter_1;
input 	always01;
output 	wait_latency_counter_0;
output 	mem_used_1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	entries_1;
input 	entries_0;
input 	d_read;
output 	nios2_data_master_waitrequest;
output 	av_begintransfer;
output 	sink_ready;
output 	saved_grant_0;
output 	WideOr0;
output 	saved_grant_01;
output 	mem_used_11;
output 	Equal5;
output 	saved_grant_02;
input 	waitrequest;
output 	mem_used_12;
input 	av_waitrequest;
output 	mem_used_13;
output 	WideOr01;
output 	src0_valid;
input 	za_valid;
output 	src0_valid1;
output 	read_latency_shift_reg_0;
output 	WideOr1;
output 	WideOr11;
output 	av_waitrequest1;
output 	Equal1;
output 	src5_valid;
output 	saved_grant_1;
input 	i_read;
input 	F_pc_25;
output 	src_valid;
output 	src_data_68;
output 	src_data_58;
output 	src_valid1;
output 	src_data_59;
output 	src_data_60;
output 	src_data_61;
output 	src_data_48;
output 	src_data_62;
output 	src_data_49;
output 	src_data_50;
output 	src_data_51;
output 	m0_write;
output 	m0_write1;
output 	src_data_52;
output 	src_data_53;
output 	src_data_54;
output 	src_data_55;
output 	src_data_56;
output 	src_data_57;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	src_valid2;
output 	rf_source_valid;
output 	read_latency_shift_reg;
output 	src1_valid;
output 	src1_valid1;
output 	src1_valid2;
output 	WideOr12;
input 	hbreak_enabled;
output 	src0_valid2;
output 	av_readdata_pre_0;
input 	za_data_0;
input 	address_reg_a_0;
output 	src_data_0;
output 	av_readdata_pre_221;
output 	av_readdata_pre_23;
input 	za_data_24;
output 	av_readdata_pre_24;
input 	za_data_25;
output 	av_readdata_pre_25;
input 	za_data_26;
output 	av_readdata_pre_26;
input 	za_data_1;
output 	av_readdata_pre_1;
input 	za_data_4;
output 	av_readdata_pre_4;
input 	za_data_3;
output 	av_readdata_pre_3;
input 	za_data_2;
output 	av_readdata_pre_2;
output 	WideOr13;
output 	src_data_461;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_161;
input 	za_data_5;
output 	av_readdata_pre_5;
output 	av_readdata_pre_8;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
input 	za_data_28;
output 	av_readdata_pre_28;
output 	av_readdata_pre_211;
input 	za_data_29;
output 	av_readdata_pre_29;
input 	za_data_30;
output 	av_readdata_pre_30;
input 	za_data_31;
output 	av_readdata_pre_31;
output 	av_readdata_pre_171;
output 	av_readdata_pre_181;
input 	za_data_27;
output 	av_readdata_pre_27;
input 	za_data_7;
output 	av_readdata_pre_7;
input 	za_data_6;
output 	av_readdata_pre_6;
output 	av_readdata_pre_201;
output 	av_readdata_pre_191;
output 	src_data_1;
output 	src_data_2;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
output 	src_data_6;
output 	src_data_7;
input 	b_full;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
input 	d_writedata_24;
output 	src_payload24;
input 	d_writedata_25;
output 	src_payload25;
input 	d_writedata_26;
output 	src_payload26;
input 	d_writedata_27;
output 	src_payload27;
input 	d_writedata_28;
output 	src_payload28;
input 	d_writedata_29;
output 	src_payload29;
input 	d_writedata_30;
output 	src_payload30;
input 	d_writedata_31;
output 	src_payload31;
input 	readdata_01;
output 	src_data_511;
output 	src_payload32;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_462;
output 	src_data_471;
output 	src_data_481;
output 	src_data_491;
output 	src_data_501;
output 	src_data_32;
input 	ien_AF;
input 	read_0;
input 	readdata_02;
output 	av_readdata_pre_81;
input 	ien_AE;
input 	av_readdata_9;
input 	av_readdata_8;
output 	src_payload33;
output 	src_data_34;
output 	src_payload34;
output 	src_payload35;
output 	src_data_35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_data_33;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_payload48;
output 	src_payload49;
output 	src_payload50;
output 	src_payload51;
output 	av_readdata_pre_91;
output 	src_payload52;
output 	src_data_24;
output 	src_payload53;
output 	src_payload54;
output 	src_data_25;
output 	src_payload55;
output 	src_data_26;
output 	src_payload56;
output 	src_data_27;
output 	src_payload57;
output 	src_data_28;
output 	src_payload58;
output 	src_payload59;
output 	src_payload60;
output 	src_payload61;
output 	src_payload62;
output 	av_readdata_pre_151;
output 	src_payload63;
output 	av_readdata_pre_141;
output 	av_readdata_pre_131;
output 	av_readdata_pre_121;
output 	av_readdata_pre_101;
input 	readdata_110;
input 	readdata_111;
input 	readdata_210;
input 	readdata_211;
input 	readdata_32;
input 	readdata_33;
input 	readdata_41;
input 	readdata_42;
input 	readdata_51;
input 	readdata_52;
input 	readdata_61;
input 	readdata_62;
input 	readdata_71;
input 	readdata_72;
input 	b_non_empty;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
output 	src_payload64;
output 	src_data_382;
output 	src_data_402;
output 	src_data_392;
output 	src_data_452;
output 	src_data_442;
output 	src_data_432;
output 	src_data_422;
output 	src_data_412;
output 	src_payload65;
output 	src_data_321;
input 	b_full1;
output 	src_data_29;
output 	src_data_30;
output 	src_data_31;
input 	rvalid;
input 	woverflow;
input 	ac;
output 	src_payload66;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_data_341;
output 	src_payload70;
output 	src_payload71;
output 	src_data_351;
output 	src_payload72;
output 	src_payload73;
output 	src_payload74;
output 	src_payload75;
output 	src_data_331;
output 	src_payload76;
output 	src_payload77;
output 	src_payload78;
output 	src_payload79;
output 	src_payload80;
output 	src_payload81;
output 	src_payload82;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_payload86;
output 	src_payload87;
output 	src_payload88;
output 	src_payload89;
output 	src_payload90;
output 	src_payload91;
output 	src_payload92;
output 	src_payload93;
output 	src_payload94;
output 	src_payload95;
output 	src_payload96;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \router|Equal1~0_combout ;
wire \router|Equal1~1_combout ;
wire \router|Equal2~0_combout ;
wire \sw_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \sw_s1_translator|wait_latency_counter[1]~q ;
wire \sw_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_data_master_translator|read_accepted~q ;
wire \router|always1~0_combout ;
wire \sw_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \led_s1_agent|m0_write~0_combout ;
wire \led_s1_translator|read_latency_shift_reg~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem_used[7]~q ;
wire \router|Equal1~2_combout ;
wire \router|Equal2~1_combout ;
wire \cmd_demux|src5_valid~0_combout ;
wire \nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \ram_s1_translator|read_latency_shift_reg[0]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][86]~q ;
wire \ram_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][86]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \led_s1_translator|read_latency_shift_reg[0]~q ;
wire \sw_s1_translator|read_latency_shift_reg[0]~q ;
wire \nios2_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \nios2_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \nios2_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \led_s1_agent|m0_write~1_combout ;
wire \nios2_data_master_translator|uav_read~0_combout ;
wire \nios2_instruction_master_translator|read_accepted~q ;
wire \nios2_instruction_master_agent|cp_valid~0_combout ;
wire \router_001|Equal1~0_combout ;
wire \router_001|Equal1~1_combout ;
wire \router_001|Equal1~2_combout ;
wire \router_001|Equal2~0_combout ;
wire \router_001|Equal2~1_combout ;
wire \sw_s1_agent|m0_write~1_combout ;
wire \sw_s1_translator|av_waitrequest_generated~0_combout ;
wire \cmd_demux_001|src2_valid~0_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \cmd_mux_004|saved_grant[1]~q ;
wire \cmd_demux|src4_valid~0_combout ;
wire \ram_s1_agent_rsp_fifo|mem~0_combout ;
wire \cmd_demux|src1_valid~0_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \nios2_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \ram_s1_translator|read_latency_shift_reg~0_combout ;
wire \router_001|Equal1~3_combout ;
wire \ram_s1_agent_rsp_fifo|mem~3_combout ;
wire \sw_s1_translator|av_readdata_pre[0]~q ;
wire \led_s1_translator|av_readdata_pre[0]~q ;
wire \cmd_demux|src5_valid~2_combout ;
wire \sw_s1_translator|av_readdata_pre[1]~q ;
wire \led_s1_translator|av_readdata_pre[1]~q ;
wire \sw_s1_translator|av_readdata_pre[2]~q ;
wire \led_s1_translator|av_readdata_pre[2]~q ;
wire \sw_s1_translator|av_readdata_pre[3]~q ;
wire \led_s1_translator|av_readdata_pre[3]~q ;
wire \sw_s1_translator|av_readdata_pre[4]~q ;
wire \led_s1_translator|av_readdata_pre[4]~q ;
wire \sw_s1_translator|av_readdata_pre[5]~q ;
wire \led_s1_translator|av_readdata_pre[5]~q ;
wire \sw_s1_translator|av_readdata_pre[6]~q ;
wire \led_s1_translator|av_readdata_pre[6]~q ;
wire \sw_s1_translator|av_readdata_pre[7]~q ;
wire \led_s1_translator|av_readdata_pre[7]~q ;


sdram_demo_sdram_demo_mm_interconnect_0_router_001 router_001(
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_18(F_pc_18),
	.F_pc_19(F_pc_19),
	.F_pc_20(F_pc_20),
	.F_pc_21(F_pc_21),
	.F_pc_22(F_pc_22),
	.F_pc_23(F_pc_23),
	.F_pc_24(F_pc_24),
	.F_pc_26(F_pc_26),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_9(F_pc_9),
	.F_pc_11(F_pc_11),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_10(F_pc_10),
	.F_pc_25(F_pc_25),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.Equal12(\router_001|Equal1~2_combout ),
	.Equal2(\router_001|Equal2~0_combout ),
	.Equal21(\router_001|Equal2~1_combout ),
	.Equal13(\router_001|Equal1~3_combout ));

sdram_demo_sdram_demo_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.src1_valid(src1_valid),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.WideOr1(WideOr12));

sdram_demo_sdram_demo_mm_interconnect_0_rsp_mux rsp_mux(
	.ram_block1a32(ram_block1a32),
	.ram_block1a0(ram_block1a0),
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.ram_block1a56(ram_block1a56),
	.ram_block1a24(ram_block1a24),
	.ram_block1a57(ram_block1a57),
	.ram_block1a25(ram_block1a25),
	.ram_block1a58(ram_block1a58),
	.ram_block1a26(ram_block1a26),
	.ram_block1a33(ram_block1a33),
	.ram_block1a1(ram_block1a1),
	.ram_block1a36(ram_block1a36),
	.ram_block1a4(ram_block1a4),
	.ram_block1a35(ram_block1a35),
	.ram_block1a3(ram_block1a3),
	.ram_block1a34(ram_block1a34),
	.ram_block1a2(ram_block1a2),
	.ram_block1a37(ram_block1a37),
	.ram_block1a5(ram_block1a5),
	.ram_block1a60(ram_block1a60),
	.ram_block1a28(ram_block1a28),
	.ram_block1a61(ram_block1a61),
	.ram_block1a29(ram_block1a29),
	.ram_block1a62(ram_block1a62),
	.ram_block1a30(ram_block1a30),
	.ram_block1a63(ram_block1a63),
	.ram_block1a31(ram_block1a31),
	.ram_block1a59(ram_block1a59),
	.ram_block1a27(ram_block1a27),
	.ram_block1a39(ram_block1a39),
	.ram_block1a7(ram_block1a7),
	.ram_block1a38(ram_block1a38),
	.ram_block1a6(ram_block1a6),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(read_latency_shift_reg_0),
	.read_latency_shift_reg_02(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\nios2_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.WideOr11(WideOr1),
	.WideOr12(WideOr11),
	.src0_valid2(src0_valid2),
	.av_readdata_pre_01(av_readdata_pre_0),
	.za_data_0(za_data_0),
	.av_readdata_pre_02(\sw_s1_translator|av_readdata_pre[0]~q ),
	.address_reg_a_0(address_reg_a_0),
	.av_readdata_pre_03(\led_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.za_data_24(za_data_24),
	.av_readdata_pre_24(av_readdata_pre_24),
	.za_data_25(za_data_25),
	.av_readdata_pre_25(av_readdata_pre_25),
	.za_data_26(za_data_26),
	.av_readdata_pre_26(av_readdata_pre_26),
	.za_data_1(za_data_1),
	.av_readdata_pre_11(av_readdata_pre_1),
	.za_data_4(za_data_4),
	.av_readdata_pre_41(av_readdata_pre_4),
	.za_data_3(za_data_3),
	.av_readdata_pre_31(av_readdata_pre_3),
	.za_data_2(za_data_2),
	.av_readdata_pre_21(av_readdata_pre_2),
	.za_data_5(za_data_5),
	.av_readdata_pre_51(av_readdata_pre_5),
	.za_data_28(za_data_28),
	.av_readdata_pre_28(av_readdata_pre_28),
	.za_data_29(za_data_29),
	.av_readdata_pre_29(av_readdata_pre_29),
	.za_data_30(za_data_30),
	.av_readdata_pre_30(av_readdata_pre_30),
	.za_data_31(za_data_31),
	.av_readdata_pre_311(av_readdata_pre_31),
	.za_data_27(za_data_27),
	.av_readdata_pre_27(av_readdata_pre_27),
	.za_data_7(za_data_7),
	.av_readdata_pre_71(av_readdata_pre_7),
	.za_data_6(za_data_6),
	.av_readdata_pre_61(av_readdata_pre_6),
	.av_readdata_pre_12(\sw_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_13(\led_s1_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_22(\sw_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_23(\led_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_32(\sw_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\led_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_42(\sw_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\led_s1_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_52(\sw_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\led_s1_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_62(\sw_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\led_s1_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_72(\sw_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\led_s1_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.src_data_24(src_data_24),
	.src_data_25(src_data_25),
	.src_data_26(src_data_26),
	.src_data_27(src_data_27),
	.src_data_28(src_data_28),
	.src_data_29(src_data_29),
	.src_data_30(src_data_30),
	.src_data_31(src_data_31));

sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001_2 rsp_demux_005(
	.za_valid(za_valid),
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid2));

sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001_1 rsp_demux_004(
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\ram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\ram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid1));

sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001 rsp_demux_001(
	.read_latency_shift_reg_0(\nios2_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src1_valid(src1_valid),
	.src0_valid(src0_valid2));

sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001_2 cmd_mux_005(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_18(F_pc_18),
	.F_pc_19(F_pc_19),
	.F_pc_20(F_pc_20),
	.F_pc_21(F_pc_21),
	.F_pc_22(F_pc_22),
	.F_pc_23(F_pc_23),
	.F_pc_24(F_pc_24),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_9(F_pc_9),
	.F_pc_11(F_pc_11),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_10(F_pc_10),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.F_pc_8(F_pc_8),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_read(d_read),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.av_begintransfer(av_begintransfer),
	.saved_grant_0(saved_grant_0),
	.WideOr0(WideOr0),
	.src5_valid(\cmd_demux|src5_valid~0_combout ),
	.Equal1(Equal1),
	.src5_valid1(src5_valid),
	.saved_grant_1(saved_grant_1),
	.i_read(i_read),
	.read_accepted1(\nios2_instruction_master_translator|read_accepted~q ),
	.cp_valid(\nios2_instruction_master_agent|cp_valid~0_combout ),
	.Equal11(\router_001|Equal1~0_combout ),
	.Equal12(\router_001|Equal1~1_combout ),
	.Equal13(\router_001|Equal1~2_combout ),
	.Equal2(\router_001|Equal2~1_combout ),
	.src_valid(src_valid),
	.src_data_68(src_data_68),
	.src_data_58(src_data_58),
	.src_valid1(src_valid1),
	.src_data_59(src_data_59),
	.src_data_60(src_data_60),
	.src_data_61(src_data_61),
	.src_data_48(src_data_48),
	.src_data_62(src_data_62),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.src_data_51(src_data_51),
	.src_data_52(src_data_52),
	.src_data_53(src_data_53),
	.src_data_54(src_data_54),
	.src_data_55(src_data_55),
	.src_data_56(src_data_56),
	.src_data_57(src_data_57),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.src5_valid2(\cmd_demux|src5_valid~2_combout ),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.d_writedata_24(d_writedata_24),
	.src_payload24(src_payload24),
	.d_writedata_25(d_writedata_25),
	.src_payload25(src_payload25),
	.d_writedata_26(d_writedata_26),
	.src_payload26(src_payload26),
	.d_writedata_27(d_writedata_27),
	.src_payload27(src_payload27),
	.d_writedata_28(d_writedata_28),
	.src_payload28(src_payload28),
	.d_writedata_29(d_writedata_29),
	.src_payload29(src_payload29),
	.d_writedata_30(d_writedata_30),
	.src_payload30(src_payload30),
	.d_writedata_31(d_writedata_31),
	.src_payload31(src_payload31),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001_1 cmd_mux_004(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.F_pc_9(F_pc_9),
	.F_pc_11(F_pc_11),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_10(F_pc_10),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.F_pc_8(F_pc_8),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_11),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.cp_valid(\nios2_instruction_master_agent|cp_valid~0_combout ),
	.Equal11(\router_001|Equal1~0_combout ),
	.Equal12(\router_001|Equal1~1_combout ),
	.Equal13(\router_001|Equal1~2_combout ),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.src_valid(src_valid2),
	.src4_valid(\cmd_demux|src4_valid~0_combout ),
	.read_latency_shift_reg(\ram_s1_translator|read_latency_shift_reg~0_combout ),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.src_data_51(src_data_511),
	.src_payload(src_payload32),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_46(src_data_462),
	.src_data_47(src_data_471),
	.src_data_48(src_data_481),
	.src_data_49(src_data_491),
	.src_data_50(src_data_501),
	.src_data_32(src_data_32),
	.src_payload1(src_payload33),
	.src_data_34(src_data_34),
	.src_payload2(src_payload34),
	.src_payload3(src_payload35),
	.src_data_35(src_data_35),
	.src_payload4(src_payload36),
	.src_payload5(src_payload37),
	.src_payload6(src_payload38),
	.src_payload7(src_payload39),
	.src_payload8(src_payload40),
	.src_payload9(src_payload41),
	.src_payload10(src_payload42),
	.src_data_33(src_data_33),
	.src_payload11(src_payload43),
	.src_payload12(src_payload44),
	.src_payload13(src_payload45),
	.src_payload14(src_payload46),
	.src_payload15(src_payload47),
	.src_payload16(src_payload48),
	.src_payload17(src_payload49),
	.src_payload18(src_payload50),
	.src_payload19(src_payload51),
	.src_payload20(src_payload52),
	.src_payload21(src_payload53),
	.src_payload22(src_payload54),
	.src_payload23(src_payload55),
	.src_payload24(src_payload56),
	.src_payload25(src_payload57),
	.src_payload26(src_payload58),
	.src_payload27(src_payload59),
	.src_payload28(src_payload60),
	.src_payload29(src_payload61),
	.src_payload30(src_payload62),
	.src_payload31(src_payload63),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001 cmd_mux_001(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.F_pc_8(F_pc_8),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.saved_grant_0(saved_grant_02),
	.write(\nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.hbreak_enabled(hbreak_enabled),
	.WideOr11(WideOr13),
	.src_data_46(src_data_461),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.src_payload(src_payload64),
	.src_data_38(src_data_382),
	.src_data_40(src_data_402),
	.src_data_39(src_data_392),
	.src_data_45(src_data_452),
	.src_data_44(src_data_442),
	.src_data_43(src_data_432),
	.src_data_42(src_data_422),
	.src_data_41(src_data_412),
	.src_payload1(src_payload65),
	.src_data_32(src_data_321),
	.src_payload2(src_payload66),
	.src_payload3(src_payload67),
	.src_payload4(src_payload68),
	.src_payload5(src_payload69),
	.src_data_34(src_data_341),
	.src_payload6(src_payload70),
	.src_payload7(src_payload71),
	.src_data_35(src_data_351),
	.src_payload8(src_payload72),
	.src_payload9(src_payload73),
	.src_payload10(src_payload74),
	.src_payload11(src_payload75),
	.src_data_33(src_data_331),
	.src_payload12(src_payload76),
	.src_payload13(src_payload77),
	.src_payload14(src_payload78),
	.src_payload15(src_payload79),
	.src_payload16(src_payload80),
	.src_payload17(src_payload81),
	.src_payload18(src_payload82),
	.src_payload19(src_payload83),
	.src_payload20(src_payload84),
	.src_payload21(src_payload85),
	.src_payload22(src_payload86),
	.src_payload23(src_payload87),
	.src_payload24(src_payload88),
	.src_payload25(src_payload89),
	.src_payload26(src_payload90),
	.src_payload27(src_payload91),
	.src_payload28(src_payload92),
	.src_payload29(src_payload93),
	.src_payload30(src_payload94),
	.src_payload31(src_payload95),
	.src_payload32(src_payload96),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.F_pc_9(F_pc_9),
	.cp_valid(\nios2_instruction_master_agent|cp_valid~0_combout ),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.Equal12(\router_001|Equal1~2_combout ),
	.Equal2(\router_001|Equal2~0_combout ),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ));

sdram_demo_sdram_demo_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.always0(always0),
	.Equal1(\router|Equal1~0_combout ),
	.Equal11(\router|Equal1~1_combout ),
	.Equal2(\router|Equal2~0_combout ),
	.Equal4(Equal4),
	.rst1(rst1),
	.mem_used_1(mem_used_1),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.d_read(d_read),
	.mem_used_11(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\sw_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sw_s1_translator|wait_latency_counter[0]~q ),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.av_begintransfer(av_begintransfer),
	.m0_write(\sw_s1_agent|m0_write~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.sink_ready1(sink_ready),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_0(saved_grant_0),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.WideOr0(WideOr0),
	.Equal12(\router|Equal1~2_combout ),
	.saved_grant_01(saved_grant_01),
	.mem_used_12(mem_used_11),
	.Equal21(\router|Equal2~1_combout ),
	.Equal5(Equal5),
	.src5_valid(\cmd_demux|src5_valid~0_combout ),
	.saved_grant_02(saved_grant_02),
	.write(\nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest(av_waitrequest),
	.mem_used_13(mem_used_13),
	.WideOr01(WideOr01),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.Equal13(Equal1),
	.src5_valid1(src5_valid),
	.src4_valid(\cmd_demux|src4_valid~0_combout ),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src5_valid2(\cmd_demux|src5_valid~2_combout ));

sdram_demo_sdram_demo_mm_interconnect_0_router router(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_3(W_alu_result_3),
	.Equal1(\router|Equal1~0_combout ),
	.Equal11(\router|Equal1~1_combout ),
	.Equal2(\router|Equal2~0_combout ),
	.Equal4(Equal4),
	.d_read(d_read),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.always1(\router|always1~0_combout ),
	.Equal12(\router|Equal1~2_combout ),
	.Equal21(\router|Equal2~1_combout ),
	.Equal5(Equal5),
	.Equal13(Equal1));

sdram_demo_altera_avalon_sc_fifo_4 sdram_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.WideOr0(WideOr0),
	.za_valid(za_valid),
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.saved_grant_1(saved_grant_1),
	.src_valid(src_valid),
	.src_data_68(src_data_68),
	.src_valid1(src_valid1),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_agent_4 sdram_s1_agent(
	.always0(always0),
	.saved_grant_0(saved_grant_0),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.m0_write(m0_write),
	.m0_write1(m0_write1));

sdram_demo_altera_avalon_sc_fifo_3 ram_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\ram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\ram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.i_read(i_read),
	.read_accepted(\nios2_instruction_master_translator|read_accepted~q ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.src_valid(src_valid2),
	.src4_valid(\cmd_demux|src4_valid~0_combout ),
	.mem(\ram_s1_agent_rsp_fifo|mem~0_combout ),
	.read_latency_shift_reg(\ram_s1_translator|read_latency_shift_reg~0_combout ),
	.mem1(\ram_s1_agent_rsp_fifo|mem~3_combout ),
	.clk(clk_clk));

sdram_demo_altera_avalon_sc_fifo_5 sw_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.read_latency_shift_reg_0(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.av_waitrequest_generated(\sw_s1_translator|av_waitrequest_generated~0_combout ),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_agent_5 sw_s1_agent(
	.Equal4(Equal4),
	.mem_used_1(\sw_s1_agent_rsp_fifo|mem_used[1]~q ),
	.av_begintransfer(av_begintransfer),
	.always1(\router|always1~0_combout ),
	.m0_write(\sw_s1_agent|m0_write~0_combout ),
	.m0_write1(\sw_s1_agent|m0_write~1_combout ));

sdram_demo_altera_avalon_sc_fifo_1 led_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.clk(clk_clk));

sdram_demo_altera_merlin_master_translator_1 nios2_instruction_master_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.WideOr0(WideOr0),
	.write(\nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(saved_grant_1),
	.i_read(i_read),
	.read_accepted1(\nios2_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~2_combout ),
	.Equal2(\router_001|Equal2~1_combout ),
	.saved_grant_11(\cmd_mux_001|saved_grant[1]~q ),
	.WideOr1(WideOr12),
	.Equal11(\router_001|Equal1~3_combout ),
	.mem(\ram_s1_agent_rsp_fifo|mem~3_combout ),
	.clk(clk_clk));

sdram_demo_altera_merlin_master_translator nios2_data_master_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted1(write_accepted),
	.always0(always0),
	.rst1(rst1),
	.d_read(d_read),
	.av_waitrequest(nios2_data_master_waitrequest),
	.read_accepted1(\nios2_data_master_translator|read_accepted~q ),
	.sink_ready(sink_ready),
	.WideOr0(WideOr01),
	.WideOr1(WideOr11),
	.av_waitrequest1(av_waitrequest1),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_translator_3 ram_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\ram_s1_translator|read_latency_shift_reg[0]~q ),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid2),
	.mem(\ram_s1_agent_rsp_fifo|mem~0_combout ),
	.read_latency_shift_reg(\ram_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_translator_5 sw_s1_translator(
	.reset(r_sync_rst),
	.always0(always0),
	.Equal4(Equal4),
	.wait_latency_counter_1(\sw_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sw_s1_translator|wait_latency_counter[0]~q ),
	.always1(\router|always1~0_combout ),
	.m0_write(\sw_s1_agent|m0_write~0_combout ),
	.sink_ready(sink_ready),
	.read_latency_shift_reg_0(\sw_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\sw_s1_agent|m0_write~1_combout ),
	.av_waitrequest_generated(\sw_s1_translator|av_waitrequest_generated~0_combout ),
	.av_readdata_pre_0(\sw_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\sw_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\sw_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\sw_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\sw_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\sw_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\sw_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\sw_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_71,readdata_61,readdata_51,readdata_41,readdata_32,readdata_210,readdata_110,readdata_01}),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_translator_1 led_s1_translator(
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.always0(always0),
	.Equal4(Equal4),
	.wait_latency_counter_1(wait_latency_counter_1),
	.always01(always01),
	.wait_latency_counter_0(wait_latency_counter_0),
	.mem_used_1(mem_used_1),
	.m0_write(\led_s1_agent|m0_write~0_combout ),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(\led_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\led_s1_agent|m0_write~1_combout ),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.av_readdata_pre_0(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\led_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\led_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\led_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\led_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\led_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\led_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\led_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_72,readdata_62,readdata_52,readdata_42,readdata_33,readdata_211,readdata_111,readdata_02}),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_translator_2 nios2_debug_mem_slave_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.rst1(rst1),
	.write(\nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.read_latency_shift_reg_0(\nios2_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.rf_source_valid(rf_source_valid),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_22(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_16(av_readdata_pre_161),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_21(av_readdata_pre_211),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_17(av_readdata_pre_171),
	.av_readdata_pre_18(av_readdata_pre_181),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_20(av_readdata_pre_201),
	.av_readdata_pre_19(av_readdata_pre_191),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_translator jtag_uart_avalon_jtag_slave_translator(
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.q_b_0(q_b_0),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_16(av_readdata_pre_16),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Add13,Add12,Add1,Add11,Add14,Add15,Add16,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,GND_port,GND_port,GND_port,GND_port,GND_port,GND_port,ien_AE,ien_AF}),
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.rst1(rst1),
	.d_read(d_read),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.av_begintransfer(av_begintransfer),
	.Equal5(Equal5),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.b_full(b_full),
	.read_0(read_0),
	.av_readdata_pre_8(av_readdata_pre_81),
	.av_readdata_pre_9(av_readdata_pre_91),
	.av_readdata_pre_15(av_readdata_pre_151),
	.av_readdata_pre_14(av_readdata_pre_141),
	.av_readdata_pre_13(av_readdata_pre_131),
	.av_readdata_pre_12(av_readdata_pre_121),
	.av_readdata_pre_10(av_readdata_pre_101),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.b_full1(b_full1),
	.clk(clk_clk));

sdram_demo_altera_merlin_master_agent_1 nios2_instruction_master_agent(
	.rst1(rst1),
	.i_read(i_read),
	.read_accepted(\nios2_instruction_master_translator|read_accepted~q ),
	.cp_valid(\nios2_instruction_master_agent|cp_valid~0_combout ));

sdram_demo_altera_merlin_slave_agent_1 led_s1_agent(
	.W_alu_result_4(W_alu_result_4),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.Equal4(Equal4),
	.rst1(rst1),
	.mem_used_1(mem_used_1),
	.d_read(d_read),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.m0_write(\led_s1_agent|m0_write~0_combout ),
	.m0_write1(\led_s1_agent|m0_write~1_combout ));

sdram_demo_altera_avalon_sc_fifo_2 nios2_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_02),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_12),
	.write(\nios2_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.read_latency_shift_reg_0(\nios2_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\nios2_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.uav_read(\nios2_data_master_translator|uav_read~0_combout ),
	.i_read(i_read),
	.read_accepted(\nios2_instruction_master_translator|read_accepted~q ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.mem(\nios2_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.rf_source_valid(rf_source_valid),
	.clk(clk_clk));

sdram_demo_altera_merlin_slave_agent_2 nios2_debug_mem_slave_agent(
	.saved_grant_0(saved_grant_02),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.mem(\nios2_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.rf_source_valid(rf_source_valid));

sdram_demo_altera_avalon_sc_fifo jtag_uart_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.d_read(d_read),
	.read_accepted(\nios2_data_master_translator|read_accepted~q ),
	.Equal5(Equal5),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.clk(clk_clk));

endmodule

module sdram_demo_altera_avalon_sc_fifo (
	reset,
	rst1,
	d_read,
	read_accepted,
	Equal5,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	d_read;
input 	read_accepted;
input 	Equal5;
input 	av_waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~0_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!rst1),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(!Equal5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!av_waitrequest),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!av_waitrequest),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hF377FFFFF377FFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_avalon_sc_fifo_1 (
	reset,
	mem_used_1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	uav_read,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	uav_read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!uav_read),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!uav_read),
	.datac(!read_latency_shift_reg_0),
	.datad(!\mem_used[0]~q ),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hF377FFFFF377FFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_avalon_sc_fifo_2 (
	reset,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	write,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	uav_read,
	i_read,
	read_accepted,
	saved_grant_1,
	mem,
	rf_source_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
output 	write;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
input 	uav_read;
input 	i_read;
input 	read_accepted;
input 	saved_grant_1;
output 	mem;
input 	rf_source_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!read_accepted),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg_0),
	.datad(!rf_source_valid),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hB8FFFFFFB8FFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg_0),
	.datad(!rf_source_valid),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBBFFF3FFBBFFF3FF;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

endmodule

module sdram_demo_altera_avalon_sc_fifo_3 (
	reset,
	rst1,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	uav_read,
	i_read,
	read_accepted,
	saved_grant_1,
	src_valid,
	src4_valid,
	mem,
	read_latency_shift_reg,
	mem1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_0;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
input 	uav_read;
input 	i_read;
input 	read_accepted;
input 	saved_grant_1;
input 	src_valid;
input 	src4_valid;
output 	mem;
input 	read_latency_shift_reg;
output 	mem1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!read_accepted),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem1),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~3 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~4 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~4 .extended_lut = "off";
defparam \mem_used[0]~4 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \mem_used[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~5 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src4_valid),
	.datad(!src_valid),
	.datae(!mem),
	.dataf(!\mem_used[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~5 .extended_lut = "off";
defparam \mem_used[0]~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[0]~5 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!rst1),
	.datab(!\mem_used[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~3 (
	.dataa(!saved_grant_0),
	.datab(!src4_valid),
	.datac(!src_valid),
	.datad(!mem),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(!\mem_used[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~3 .extended_lut = "off";
defparam \mem_used[1]~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[1]~3 .shared_arith = "off";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

endmodule

module sdram_demo_altera_avalon_sc_fifo_4 (
	reset,
	saved_grant_0,
	mem_used_7,
	WideOr0,
	za_valid,
	mem_86_0,
	mem_68_0,
	Equal1,
	src5_valid,
	saved_grant_1,
	src_valid,
	src_data_68,
	src_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
output 	mem_used_7;
input 	WideOr0;
input 	za_valid;
output 	mem_86_0;
output 	mem_68_0;
input 	Equal1;
input 	src5_valid;
input 	saved_grant_1;
input 	src_valid;
input 	src_data_68;
input 	src_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used~3_combout ;
wire \mem_used[6]~4_combout ;
wire \mem_used[6]~q ;
wire \mem_used~6_combout ;
wire \mem_used[5]~q ;
wire \mem_used~8_combout ;
wire \mem_used[4]~q ;
wire \mem_used~9_combout ;
wire \mem_used[3]~q ;
wire \mem_used~7_combout ;
wire \mem_used[2]~q ;
wire \mem_used~5_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[7]~0_combout ;
wire \mem[7][86]~q ;
wire \mem~12_combout ;
wire \always6~0_combout ;
wire \mem[6][86]~q ;
wire \mem~10_combout ;
wire \always5~0_combout ;
wire \mem[5][86]~q ;
wire \mem~8_combout ;
wire \always4~0_combout ;
wire \mem[4][86]~q ;
wire \mem~6_combout ;
wire \always3~0_combout ;
wire \mem[3][86]~q ;
wire \mem~4_combout ;
wire \always2~0_combout ;
wire \mem[2][86]~q ;
wire \mem~2_combout ;
wire \always1~0_combout ;
wire \mem[1][86]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[7][68]~q ;
wire \mem~13_combout ;
wire \mem[6][68]~q ;
wire \mem~11_combout ;
wire \mem[5][68]~q ;
wire \mem~9_combout ;
wire \mem[4][68]~q ;
wire \mem~7_combout ;
wire \mem[3][68]~q ;
wire \mem~5_combout ;
wire \mem[2][68]~q ;
wire \mem~3_combout ;
wire \mem[1][68]~q ;
wire \mem~1_combout ;


dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!saved_grant_0),
	.datab(!WideOr0),
	.datac(!Equal1),
	.datad(!src5_valid),
	.datae(!src_valid),
	.dataf(!src_data_68),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used~3 (
	.dataa(!mem_used_7),
	.datab(!WideOr0),
	.datac(!src_valid1),
	.datad(!src_valid),
	.datae(!src_data_68),
	.dataf(!\mem_used[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~3 .extended_lut = "off";
defparam \mem_used~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used~3 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[6]~4 (
	.dataa(!WideOr0),
	.datab(!za_valid),
	.datac(!src_valid1),
	.datad(!src_valid),
	.datae(!src_data_68),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[6]~4 .extended_lut = "off";
defparam \mem_used[6]~4 .lut_mask = 64'h6996966996696996;
defparam \mem_used[6]~4 .shared_arith = "off";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cyclonev_lcell_comb \mem_used~6 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[6]~q ),
	.dataf(!\mem_used[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~6 .extended_lut = "off";
defparam \mem_used~6 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \mem_used~6 .shared_arith = "off";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cyclonev_lcell_comb \mem_used~8 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[5]~q ),
	.dataf(!\mem_used[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~8 .extended_lut = "off";
defparam \mem_used~8 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \mem_used~8 .shared_arith = "off";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cyclonev_lcell_comb \mem_used~9 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[2]~q ),
	.dataf(!\mem_used[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~9 .extended_lut = "off";
defparam \mem_used~9 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \mem_used~9 .shared_arith = "off";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cyclonev_lcell_comb \mem_used~7 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[1]~q ),
	.dataf(!\mem_used[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~7 .extended_lut = "off";
defparam \mem_used~7 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \mem_used~7 .shared_arith = "off";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cyclonev_lcell_comb \mem_used~5 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[0]~q ),
	.dataf(!\mem_used[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~5 .extended_lut = "off";
defparam \mem_used~5 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \mem_used~5 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~4_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \mem_used[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!src_data_68),
	.datae(!\mem_used[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[7]~0 (
	.dataa(!mem_used_7),
	.datab(!za_valid),
	.datac(!\write~0_combout ),
	.datad(!\mem_used[0]~q ),
	.datae(!\mem_used[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[7]~0 .extended_lut = "off";
defparam \mem_used[7]~0 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \mem_used[7]~0 .shared_arith = "off";

dffeas \mem[7][86] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][86]~q ),
	.prn(vcc));
defparam \mem[7][86] .is_wysiwyg = "true";
defparam \mem[7][86] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_7),
	.datab(!saved_grant_1),
	.datac(!\mem[7][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h2727272727272727;
defparam \mem~12 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always6~0 .shared_arith = "off";

dffeas \mem[6][86] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][86]~q ),
	.prn(vcc));
defparam \mem[6][86] .is_wysiwyg = "true";
defparam \mem[6][86] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!saved_grant_1),
	.datab(!\mem_used[6]~q ),
	.datac(!\mem[6][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

cyclonev_lcell_comb \always5~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always5~0 .shared_arith = "off";

dffeas \mem[5][86] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][86]~q ),
	.prn(vcc));
defparam \mem[5][86] .is_wysiwyg = "true";
defparam \mem[5][86] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!saved_grant_1),
	.datab(!\mem_used[5]~q ),
	.datac(!\mem[5][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

cyclonev_lcell_comb \always4~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[4][86] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][86]~q ),
	.prn(vcc));
defparam \mem[4][86] .is_wysiwyg = "true";
defparam \mem[4][86] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!saved_grant_1),
	.datab(!\mem_used[4]~q ),
	.datac(!\mem[4][86]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

cyclonev_lcell_comb \always3~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always3~0 .shared_arith = "off";

dffeas \mem[3][86] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][86]~q ),
	.prn(vcc));
defparam \mem[3][86] .is_wysiwyg = "true";
defparam \mem[3][86] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!saved_grant_1),
	.datab(!\mem[3][86]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h5353535353535353;
defparam \mem~4 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always2~0 .shared_arith = "off";

dffeas \mem[2][86] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][86]~q ),
	.prn(vcc));
defparam \mem[2][86] .is_wysiwyg = "true";
defparam \mem[2][86] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_1),
	.datab(!\mem[2][86]~q ),
	.datac(!\mem_used[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h5353535353535353;
defparam \mem~2 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always1~0 .shared_arith = "off";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!saved_grant_1),
	.datab(!\mem[1][86]~q ),
	.datac(!\mem_used[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h5353535353535353;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!za_valid),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[7][68] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][68]~q ),
	.prn(vcc));
defparam \mem[7][68] .is_wysiwyg = "true";
defparam \mem[7][68] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_7),
	.datab(!src_data_68),
	.datac(!\mem[7][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h2727272727272727;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[6][68] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][68]~q ),
	.prn(vcc));
defparam \mem[6][68] .is_wysiwyg = "true";
defparam \mem[6][68] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!src_data_68),
	.datab(!\mem_used[6]~q ),
	.datac(!\mem[6][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[5][68] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][68]~q ),
	.prn(vcc));
defparam \mem[5][68] .is_wysiwyg = "true";
defparam \mem[5][68] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!src_data_68),
	.datab(!\mem_used[5]~q ),
	.datac(!\mem[5][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[4][68] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][68]~q ),
	.prn(vcc));
defparam \mem[4][68] .is_wysiwyg = "true";
defparam \mem[4][68] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!src_data_68),
	.datab(!\mem_used[4]~q ),
	.datac(!\mem[4][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[3][68] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][68]~q ),
	.prn(vcc));
defparam \mem[3][68] .is_wysiwyg = "true";
defparam \mem[3][68] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!src_data_68),
	.datab(!\mem_used[3]~q ),
	.datac(!\mem[3][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[2][68] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][68]~q ),
	.prn(vcc));
defparam \mem[2][68] .is_wysiwyg = "true";
defparam \mem[2][68] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!src_data_68),
	.datab(!\mem_used[2]~q ),
	.datac(!\mem[2][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!src_data_68),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_avalon_sc_fifo_5 (
	reset,
	mem_used_1,
	sink_ready,
	read_latency_shift_reg_0,
	av_waitrequest_generated,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	sink_ready;
input 	read_latency_shift_reg_0;
input 	av_waitrequest_generated;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!av_waitrequest_generated),
	.datac(!sink_ready),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBF1FFFFFBF1FFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!av_waitrequest_generated),
	.datac(!sink_ready),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_master_agent_1 (
	rst1,
	i_read,
	read_accepted,
	cp_valid)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	i_read;
input 	read_accepted;
output 	cp_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \cp_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_valid~0 .extended_lut = "off";
defparam \cp_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \cp_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_master_translator (
	reset,
	d_write,
	write_accepted1,
	always0,
	rst1,
	d_read,
	av_waitrequest,
	read_accepted1,
	sink_ready,
	WideOr0,
	WideOr1,
	av_waitrequest1,
	uav_read,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
output 	write_accepted1;
input 	always0;
input 	rst1;
input 	d_read;
output 	av_waitrequest;
output 	read_accepted1;
input 	sink_ready;
input 	WideOr0;
input 	WideOr1;
output 	av_waitrequest1;
output 	uav_read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write_accepted~0_combout ;
wire \read_accepted~0_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;


dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!write_accepted1),
	.datab(!d_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \av_waitrequest~0 .shared_arith = "off";

dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!d_write),
	.datab(!write_accepted1),
	.datac(!rst1),
	.datad(!d_read),
	.datae(!\end_begintransfer~q ),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'hFF7FFFFF3F7FFFFF;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \uav_read~0 (
	.dataa(!d_read),
	.datab(!read_accepted1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(uav_read),
	.sumout(),
	.cout(),
	.shareout());
defparam \uav_read~0 .extended_lut = "off";
defparam \uav_read~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \uav_read~0 .shared_arith = "off";

cyclonev_lcell_comb \write_accepted~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!write_accepted1),
	.datad(!av_waitrequest1),
	.datae(!WideOr0),
	.dataf(!sink_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_accepted~0 .extended_lut = "off";
defparam \write_accepted~0 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \write_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!rst1),
	.datab(!d_read),
	.datac(!read_accepted1),
	.datad(!sink_ready),
	.datae(!WideOr0),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \read_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \end_begintransfer~0 (
	.dataa(!always0),
	.datab(!rst1),
	.datac(!uav_read),
	.datad(!\end_begintransfer~q ),
	.datae(!sink_ready),
	.dataf(!WideOr0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\end_begintransfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \end_begintransfer~0 .extended_lut = "off";
defparam \end_begintransfer~0 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \end_begintransfer~0 .shared_arith = "off";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

endmodule

module sdram_demo_altera_merlin_master_translator_1 (
	reset,
	rst1,
	WideOr0,
	write,
	saved_grant_1,
	i_read,
	read_accepted1,
	Equal1,
	Equal2,
	saved_grant_11,
	WideOr1,
	Equal11,
	mem,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	WideOr0;
input 	write;
input 	saved_grant_1;
input 	i_read;
output 	read_accepted1;
input 	Equal1;
input 	Equal2;
input 	saved_grant_11;
input 	WideOr1;
input 	Equal11;
input 	mem;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;
wire \read_accepted~3_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!write),
	.datab(!saved_grant_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'h7777777777777777;
defparam \read_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~1 (
	.dataa(!WideOr0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~1 .extended_lut = "off";
defparam \read_accepted~1 .lut_mask = 64'h7777777777777777;
defparam \read_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~2 (
	.dataa(!Equal11),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!mem),
	.datae(!\read_accepted~0_combout ),
	.dataf(!\read_accepted~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~2 .extended_lut = "off";
defparam \read_accepted~2 .lut_mask = 64'hFFFFFFFFFFFFFF96;
defparam \read_accepted~2 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~3 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted1),
	.datad(!WideOr1),
	.datae(!\read_accepted~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~3 .extended_lut = "off";
defparam \read_accepted~3 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \read_accepted~3 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_agent_1 (
	W_alu_result_4,
	d_write,
	write_accepted,
	Equal4,
	rst1,
	mem_used_1,
	d_read,
	read_accepted,
	m0_write,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	d_write;
input 	write_accepted;
input 	Equal4;
input 	rst1;
input 	mem_used_1;
input 	d_read;
input 	read_accepted;
output 	m0_write;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!d_write),
	.datac(!write_accepted),
	.datad(!rst1),
	.datae(!d_read),
	.dataf(!read_accepted),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFFFFFFFFFBFFFFFF;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!W_alu_result_4),
	.datab(!Equal4),
	.datac(!m0_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_agent_2 (
	saved_grant_0,
	src1_valid,
	src0_valid,
	saved_grant_1,
	mem,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_0;
input 	src1_valid;
input 	src0_valid;
input 	saved_grant_1;
input 	mem;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!saved_grant_0),
	.datab(!src1_valid),
	.datac(!src0_valid),
	.datad(!saved_grant_1),
	.datae(!mem),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_agent_4 (
	always0,
	saved_grant_0,
	mem_used_7,
	Equal1,
	src5_valid,
	src_valid,
	m0_write,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	always0;
input 	saved_grant_0;
input 	mem_used_7;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
output 	m0_write;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!always0),
	.datab(!saved_grant_0),
	.datac(!mem_used_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!saved_grant_0),
	.datab(!Equal1),
	.datac(!src5_valid),
	.datad(!src_valid),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'hFFFFFFFBFFFFFFFB;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_agent_5 (
	Equal4,
	mem_used_1,
	av_begintransfer,
	always1,
	m0_write,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	Equal4;
input 	mem_used_1;
input 	av_begintransfer;
input 	always1;
output 	m0_write;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!Equal4),
	.datab(!av_begintransfer),
	.datac(!mem_used_1),
	.datad(!always1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!av_begintransfer),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_translator (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	q_b_0,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_16,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	av_readdata,
	reset,
	d_write,
	write_accepted,
	rst1,
	d_read,
	read_accepted,
	av_begintransfer,
	Equal5,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	b_full,
	read_0,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_15,
	av_readdata_pre_14,
	av_readdata_pre_13,
	av_readdata_pre_12,
	av_readdata_pre_10,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	b_full1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	q_b_0;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_16;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	[31:0] av_readdata;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	d_read;
input 	read_accepted;
output 	av_begintransfer;
input 	Equal5;
input 	av_waitrequest;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	b_full;
input 	read_0;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_15;
output 	av_readdata_pre_14;
output 	av_readdata_pre_13;
output 	av_readdata_pre_12;
output 	av_readdata_pre_10;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	b_full1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;
wire \av_readdata_pre[13]~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(q_b_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(q_b_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_6),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(q_b_7),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

cyclonev_lcell_comb \av_begintransfer~0 (
	.dataa(!d_write),
	.datab(!write_accepted),
	.datac(!rst1),
	.datad(!d_read),
	.datae(!read_accepted),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_begintransfer),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_begintransfer~0 .extended_lut = "off";
defparam \av_begintransfer~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \av_begintransfer~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!Equal5),
	.datab(!av_waitrequest),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \av_readdata_pre[13]~0 (
	.dataa(!b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_readdata_pre[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata_pre[13]~0 .extended_lut = "off";
defparam \av_readdata_pre[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \av_readdata_pre[13]~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_translator_1 (
	W_alu_result_4,
	reset,
	always0,
	Equal4,
	wait_latency_counter_1,
	always01,
	wait_latency_counter_0,
	mem_used_1,
	m0_write,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	m0_write1,
	uav_read,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	reset;
input 	always0;
input 	Equal4;
output 	wait_latency_counter_1;
input 	always01;
output 	wait_latency_counter_0;
input 	mem_used_1;
input 	m0_write;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	m0_write1;
input 	uav_read;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!always0),
	.datac(!W_alu_result_4),
	.datad(!Equal4),
	.datae(!m0_write),
	.dataf(!always01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h9FFF6FFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!always0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!always0),
	.datac(!wait_latency_counter_1),
	.datad(!m0_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!mem_used_1),
	.datab(!uav_read),
	.datac(!read_latency_shift_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_translator_2 (
	av_readdata,
	reset,
	rst1,
	write,
	read_latency_shift_reg_0,
	rf_source_valid,
	av_readdata_pre_0,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_1,
	av_readdata_pre_4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_5,
	av_readdata_pre_8,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_28,
	av_readdata_pre_21,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_27,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_20,
	av_readdata_pre_19,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	rst1;
input 	write;
output 	read_latency_shift_reg_0;
input 	rf_source_valid;
output 	av_readdata_pre_0;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_1;
output 	av_readdata_pre_4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_5;
output 	av_readdata_pre_8;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_28;
output 	av_readdata_pre_21;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_27;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!write),
	.datac(!rf_source_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_translator_3 (
	reset,
	rst1,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	Equal1,
	src5_valid,
	src_valid,
	mem,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_0;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
input 	mem;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!Equal1),
	.datad(!src5_valid),
	.datae(!src_valid),
	.dataf(!mem),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_slave_translator_5 (
	reset,
	always0,
	Equal4,
	wait_latency_counter_1,
	wait_latency_counter_0,
	always1,
	m0_write,
	sink_ready,
	read_latency_shift_reg_0,
	m0_write1,
	av_waitrequest_generated,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	always0;
input 	Equal4;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	always1;
input 	m0_write;
input 	sink_ready;
output 	read_latency_shift_reg_0;
input 	m0_write1;
output 	av_waitrequest_generated;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!always0),
	.datab(!Equal4),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!always1),
	.dataf(!m0_write1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hF9F6F6F9F6F9F9F6;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!always0),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7DFF7DFF7DFF7DFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write),
	.datac(!av_waitrequest_generated),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_cmd_demux (
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_11,
	always0,
	Equal1,
	Equal11,
	Equal2,
	Equal4,
	rst1,
	mem_used_1,
	entries_1,
	entries_0,
	d_read,
	mem_used_11,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_accepted,
	av_begintransfer,
	m0_write,
	sink_ready,
	sink_ready1,
	read_latency_shift_reg,
	saved_grant_0,
	mem_used_7,
	WideOr0,
	Equal12,
	saved_grant_01,
	mem_used_12,
	Equal21,
	Equal5,
	src5_valid,
	saved_grant_02,
	write,
	av_waitrequest,
	mem_used_13,
	WideOr01,
	uav_read,
	Equal13,
	src5_valid1,
	src4_valid,
	src1_valid,
	src5_valid2)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	always0;
input 	Equal1;
input 	Equal11;
input 	Equal2;
input 	Equal4;
input 	rst1;
input 	mem_used_1;
input 	entries_1;
input 	entries_0;
input 	d_read;
input 	mem_used_11;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	read_accepted;
input 	av_begintransfer;
input 	m0_write;
output 	sink_ready;
output 	sink_ready1;
input 	read_latency_shift_reg;
input 	saved_grant_0;
input 	mem_used_7;
output 	WideOr0;
input 	Equal12;
input 	saved_grant_01;
input 	mem_used_12;
input 	Equal21;
input 	Equal5;
output 	src5_valid;
input 	saved_grant_02;
input 	write;
input 	av_waitrequest;
input 	mem_used_13;
output 	WideOr01;
input 	uav_read;
input 	Equal13;
output 	src5_valid1;
output 	src4_valid;
output 	src1_valid;
output 	src5_valid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~3_combout ;


cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!rst1),
	.datab(!W_alu_result_4),
	.datac(!Equal4),
	.datad(!d_read),
	.datae(!read_accepted),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!always0),
	.datab(!mem_used_11),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(!sink_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hFEFDFDFEFFFFFFFF;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!entries_1),
	.datab(!entries_0),
	.datac(!mem_used_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~0 (
	.dataa(!W_alu_result_4),
	.datab(!Equal4),
	.datac(!d_read),
	.datad(!read_accepted),
	.datae(!Equal21),
	.dataf(!Equal5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~0 .extended_lut = "off";
defparam \src5_valid~0 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \src5_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg),
	.datac(!\WideOr0~2_combout ),
	.datad(!src5_valid),
	.datae(!\WideOr0~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~1 (
	.dataa(!W_alu_result_4),
	.datab(!Equal4),
	.datac(!uav_read),
	.datad(!av_begintransfer),
	.datae(!Equal21),
	.dataf(!Equal5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~1 .extended_lut = "off";
defparam \src5_valid~1 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \src5_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src4_valid~0 (
	.dataa(!av_begintransfer),
	.datab(!Equal13),
	.datac(!src5_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src4_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src4_valid~0 .extended_lut = "off";
defparam \src4_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src4_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!W_alu_result_12),
	.datab(!W_alu_result_11),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal2),
	.dataf(!av_begintransfer),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~2 (
	.dataa(!av_begintransfer),
	.datab(!Equal13),
	.datac(!src5_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~2 .extended_lut = "off";
defparam \src5_valid~2 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \src5_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!rst1),
	.datab(!saved_grant_01),
	.datac(!mem_used_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!Equal1),
	.datab(!Equal11),
	.datac(!saved_grant_0),
	.datad(!WideOr0),
	.datae(!Equal12),
	.dataf(!\WideOr0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'h9FFF6FFFFFFFFFFF;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!saved_grant_02),
	.datab(!write),
	.datac(!Equal21),
	.datad(!Equal5),
	.datae(!av_waitrequest),
	.dataf(!mem_used_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \WideOr0~3 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_cmd_demux_001 (
	F_pc_9,
	cp_valid,
	Equal1,
	Equal11,
	Equal12,
	Equal2,
	src2_valid,
	src1_valid,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	F_pc_9;
input 	cp_valid;
input 	Equal1;
input 	Equal11;
input 	Equal12;
input 	Equal2;
output 	src2_valid;
output 	src1_valid;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!cp_valid),
	.datab(!F_pc_9),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal12),
	.dataf(!Equal2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!cp_valid),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!cp_valid),
	.datab(!F_pc_9),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src0_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_0,
	write,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	src1_valid,
	src0_valid,
	saved_grant_1,
	hbreak_enabled,
	WideOr11,
	src_data_46,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	src_payload,
	src_data_38,
	src_data_40,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_41,
	src_payload1,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_33,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_9;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_8;
input 	W_alu_result_10;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
input 	F_pc_8;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	saved_grant_0;
input 	write;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
input 	src1_valid;
input 	src0_valid;
output 	saved_grant_1;
input 	hbreak_enabled;
output 	WideOr11;
output 	src_data_46;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
output 	src_payload;
output 	src_data_38;
output 	src_data_40;
output 	src_data_39;
output 	src_data_45;
output 	src_data_44;
output 	src_data_43;
output 	src_data_42;
output 	src_data_41;
output 	src_payload1;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_payload7;
output 	src_data_35;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_data_33;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


sdram_demo_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.write(write),
	.src1_valid(src1_valid),
	.src0_valid(src0_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_0),
	.datab(!src1_valid),
	.datac(!src0_valid),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!W_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!F_pc_8),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!W_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!F_pc_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!W_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!F_pc_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!W_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!F_pc_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!W_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!F_pc_7),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!W_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!F_pc_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!W_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!F_pc_5),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!W_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!F_pc_4),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!W_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!F_pc_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_0),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!d_writedata_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!d_writedata_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!d_writedata_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_2),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_3),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!d_writedata_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!d_writedata_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!d_writedata_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!d_writedata_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src1_valid),
	.datad(!src0_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	write,
	src1_valid,
	src0_valid,
	grant_0,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	write;
input 	src1_valid;
input 	src0_valid;
output 	grant_0;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src1_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src1_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src1_valid),
	.datad(!src0_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001_1 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	d_writedata_0,
	r_sync_rst,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_0,
	mem_used_1,
	Equal1,
	src5_valid,
	cp_valid,
	Equal11,
	Equal12,
	Equal13,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	src1_valid,
	saved_grant_1,
	src_valid,
	src4_valid,
	read_latency_shift_reg,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	src_data_51,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_33,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_9;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_8;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	F_pc_9;
input 	F_pc_11;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_10;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
input 	F_pc_8;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	saved_grant_0;
input 	mem_used_1;
input 	Equal1;
input 	src5_valid;
input 	cp_valid;
input 	Equal11;
input 	Equal12;
input 	Equal13;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
input 	src1_valid;
output 	saved_grant_1;
output 	src_valid;
input 	src4_valid;
input 	read_latency_shift_reg;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
output 	src_data_51;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_32;
output 	src_payload1;
output 	src_data_34;
output 	src_payload2;
output 	src_payload3;
output 	src_data_35;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_data_33;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \update_grant~1_combout ;


sdram_demo_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.src4_valid(src4_valid),
	.read_latency_shift_reg(read_latency_shift_reg),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!cp_valid),
	.datab(!Equal11),
	.datac(!Equal12),
	.datad(!Equal13),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[51] (
	.dataa(!W_alu_result_15),
	.datab(!saved_grant_0),
	.datac(!F_pc_13),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[51] .extended_lut = "off";
defparam \src_data[51] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[51] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!W_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!F_pc_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!W_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!F_pc_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!W_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!F_pc_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!W_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!F_pc_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!W_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!F_pc_4),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!W_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!F_pc_5),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!W_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!F_pc_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!W_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!F_pc_7),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!W_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!F_pc_8),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!W_alu_result_11),
	.datab(!saved_grant_0),
	.datac(!F_pc_9),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!W_alu_result_12),
	.datab(!saved_grant_0),
	.datac(!F_pc_10),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!W_alu_result_13),
	.datab(!saved_grant_0),
	.datac(!F_pc_11),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!W_alu_result_14),
	.datab(!saved_grant_0),
	.datac(!F_pc_12),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_0),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_2),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_3),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!d_writedata_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!d_writedata_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!d_writedata_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!d_writedata_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!d_writedata_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!d_writedata_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!d_writedata_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!rst1),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \update_grant~1 (
	.dataa(!saved_grant_0),
	.datab(!Equal1),
	.datac(!src5_valid),
	.datad(!\packet_in_progress~q ),
	.datae(!src_valid),
	.dataf(!\update_grant~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~1 .extended_lut = "off";
defparam \update_grant~1 .lut_mask = 64'hFF69FF96FFFFFFFF;
defparam \update_grant~1 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	Equal1,
	src5_valid,
	src1_valid,
	grant_0,
	packet_in_progress,
	saved_grant_1,
	src4_valid,
	read_latency_shift_reg,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	Equal1;
input 	src5_valid;
input 	src1_valid;
output 	grant_0;
input 	packet_in_progress;
input 	saved_grant_1;
input 	src4_valid;
input 	read_latency_shift_reg;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!Equal1),
	.datab(!src5_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!Equal1),
	.datab(!src5_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src4_valid),
	.datad(!src1_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_cmd_mux_001_2 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_24,
	W_alu_result_25,
	W_alu_result_26,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_21,
	W_alu_result_22,
	W_alu_result_23,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_17,
	F_pc_16,
	F_pc_18,
	F_pc_19,
	F_pc_20,
	F_pc_21,
	F_pc_22,
	F_pc_23,
	F_pc_24,
	F_pc_15,
	F_pc_14,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_read,
	read_accepted,
	av_begintransfer,
	saved_grant_0,
	WideOr0,
	src5_valid,
	Equal1,
	src5_valid1,
	saved_grant_1,
	i_read,
	read_accepted1,
	cp_valid,
	Equal11,
	Equal12,
	Equal13,
	Equal2,
	src_valid,
	src_data_68,
	src_data_58,
	src_valid1,
	src_data_59,
	src_data_60,
	src_data_61,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_50,
	src_data_51,
	src_data_52,
	src_data_53,
	src_data_54,
	src_data_55,
	src_data_56,
	src_data_57,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src2_valid,
	src5_valid2,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	d_writedata_24,
	src_payload24,
	d_writedata_25,
	src_payload25,
	d_writedata_26,
	src_payload26,
	d_writedata_27,
	src_payload27,
	d_writedata_28,
	src_payload28,
	d_writedata_29,
	src_payload29,
	d_writedata_30,
	src_payload30,
	d_writedata_31,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_9;
input 	W_alu_result_24;
input 	W_alu_result_25;
input 	W_alu_result_26;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_21;
input 	W_alu_result_22;
input 	W_alu_result_23;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_8;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_18;
input 	F_pc_19;
input 	F_pc_20;
input 	F_pc_21;
input 	F_pc_22;
input 	F_pc_23;
input 	F_pc_24;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_9;
input 	F_pc_11;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_10;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
input 	F_pc_8;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_read;
input 	read_accepted;
input 	av_begintransfer;
output 	saved_grant_0;
input 	WideOr0;
input 	src5_valid;
input 	Equal1;
input 	src5_valid1;
output 	saved_grant_1;
input 	i_read;
input 	read_accepted1;
input 	cp_valid;
input 	Equal11;
input 	Equal12;
input 	Equal13;
input 	Equal2;
output 	src_valid;
output 	src_data_68;
output 	src_data_58;
output 	src_valid1;
output 	src_data_59;
output 	src_data_60;
output 	src_data_61;
output 	src_data_48;
output 	src_data_62;
output 	src_data_49;
output 	src_data_50;
output 	src_data_51;
output 	src_data_52;
output 	src_data_53;
output 	src_data_54;
output 	src_data_55;
output 	src_data_56;
output 	src_data_57;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
input 	src2_valid;
input 	src5_valid2;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
input 	d_writedata_24;
output 	src_payload24;
input 	d_writedata_25;
output 	src_payload25;
input 	d_writedata_26;
output 	src_payload26;
input 	d_writedata_27;
output 	src_payload27;
input 	d_writedata_28;
output 	src_payload28;
input 	d_writedata_29;
output 	src_payload29;
input 	d_writedata_30;
output 	src_payload30;
input 	d_writedata_31;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


sdram_demo_altera_merlin_arbitrator_2 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.WideOr0(WideOr0),
	.Equal1(Equal1),
	.src5_valid(src5_valid1),
	.saved_grant_1(saved_grant_1),
	.src2_valid(src2_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src5_valid1(src5_valid2),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!cp_valid),
	.datac(!Equal11),
	.datad(!Equal12),
	.datae(!Equal13),
	.dataf(!Equal2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[68] (
	.dataa(!d_read),
	.datab(!read_accepted),
	.datac(!saved_grant_0),
	.datad(!saved_grant_1),
	.datae(!i_read),
	.dataf(!read_accepted1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[68] .extended_lut = "off";
defparam \src_data[68] .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \src_data[68] .shared_arith = "off";

cyclonev_lcell_comb \src_data[58] (
	.dataa(!W_alu_result_22),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_58),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[58] .extended_lut = "off";
defparam \src_data[58] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[58] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!av_begintransfer),
	.datab(!saved_grant_0),
	.datac(!Equal1),
	.datad(!src5_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[59] (
	.dataa(!W_alu_result_23),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_59),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[59] .extended_lut = "off";
defparam \src_data[59] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[59] .shared_arith = "off";

cyclonev_lcell_comb \src_data[60] (
	.dataa(!W_alu_result_24),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_60),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[60] .extended_lut = "off";
defparam \src_data[60] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[60] .shared_arith = "off";

cyclonev_lcell_comb \src_data[61] (
	.dataa(!W_alu_result_25),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_61),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[61] .extended_lut = "off";
defparam \src_data[61] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[61] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!W_alu_result_12),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[62] (
	.dataa(!W_alu_result_26),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_62),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[62] .extended_lut = "off";
defparam \src_data[62] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[62] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!W_alu_result_13),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!W_alu_result_14),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[51] (
	.dataa(!W_alu_result_15),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[51] .extended_lut = "off";
defparam \src_data[51] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[51] .shared_arith = "off";

cyclonev_lcell_comb \src_data[52] (
	.dataa(!W_alu_result_16),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_52),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[52] .extended_lut = "off";
defparam \src_data[52] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[52] .shared_arith = "off";

cyclonev_lcell_comb \src_data[53] (
	.dataa(!W_alu_result_17),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_53),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[53] .extended_lut = "off";
defparam \src_data[53] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[53] .shared_arith = "off";

cyclonev_lcell_comb \src_data[54] (
	.dataa(!W_alu_result_18),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_54),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[54] .extended_lut = "off";
defparam \src_data[54] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[54] .shared_arith = "off";

cyclonev_lcell_comb \src_data[55] (
	.dataa(!W_alu_result_19),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_55),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[55] .extended_lut = "off";
defparam \src_data[55] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[55] .shared_arith = "off";

cyclonev_lcell_comb \src_data[56] (
	.dataa(!W_alu_result_20),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_56),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[56] .extended_lut = "off";
defparam \src_data[56] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[56] .shared_arith = "off";

cyclonev_lcell_comb \src_data[57] (
	.dataa(!W_alu_result_21),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_57),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[57] .extended_lut = "off";
defparam \src_data[57] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[57] .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!W_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!W_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!W_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!W_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!W_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!W_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!W_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!W_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!W_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!W_alu_result_11),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!F_pc_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!d_writedata_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!d_writedata_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!d_writedata_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!d_writedata_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!d_writedata_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!d_writedata_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!d_writedata_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!WideOr0),
	.datac(!src_valid1),
	.datad(!saved_grant_1),
	.datae(!src_valid),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_merlin_arbitrator_2 (
	reset,
	saved_grant_0,
	WideOr0,
	Equal1,
	src5_valid,
	saved_grant_1,
	src2_valid,
	grant_0,
	packet_in_progress,
	grant_1,
	src5_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	WideOr0;
input 	Equal1;
input 	src5_valid;
input 	saved_grant_1;
input 	src2_valid;
output 	grant_0;
input 	packet_in_progress;
output 	grant_1;
input 	src5_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!Equal1),
	.datab(!src5_valid),
	.datac(!src2_valid),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!\top_priority_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!Equal1),
	.datab(!src5_valid),
	.datac(!src2_valid),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!\top_priority_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!WideOr0),
	.datac(!src5_valid1),
	.datad(!saved_grant_1),
	.datae(!src2_valid),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_router (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_24,
	W_alu_result_25,
	W_alu_result_26,
	W_alu_result_27,
	W_alu_result_28,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_21,
	W_alu_result_22,
	W_alu_result_23,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_3,
	Equal1,
	Equal11,
	Equal2,
	Equal4,
	d_read,
	read_accepted,
	always1,
	Equal12,
	Equal21,
	Equal5,
	Equal13)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_9;
input 	W_alu_result_24;
input 	W_alu_result_25;
input 	W_alu_result_26;
input 	W_alu_result_27;
input 	W_alu_result_28;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_21;
input 	W_alu_result_22;
input 	W_alu_result_23;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_8;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_3;
output 	Equal1;
output 	Equal11;
output 	Equal2;
output 	Equal4;
input 	d_read;
input 	read_accepted;
output 	always1;
output 	Equal12;
output 	Equal21;
output 	Equal5;
output 	Equal13;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal4~0_combout ;
wire \Equal5~0_combout ;


cyclonev_lcell_comb \Equal1~0 (
	.dataa(!W_alu_result_24),
	.datab(!W_alu_result_25),
	.datac(!W_alu_result_26),
	.datad(!W_alu_result_27),
	.datae(!W_alu_result_28),
	.dataf(!W_alu_result_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!W_alu_result_19),
	.datab(!W_alu_result_21),
	.datac(!W_alu_result_22),
	.datad(!W_alu_result_23),
	.datae(!W_alu_result_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!W_alu_result_17),
	.datab(!W_alu_result_16),
	.datac(!W_alu_result_15),
	.datad(!W_alu_result_14),
	.datae(!W_alu_result_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!W_alu_result_5),
	.datab(!W_alu_result_9),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal2),
	.dataf(!\Equal4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!W_alu_result_4),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~2 (
	.dataa(!W_alu_result_17),
	.datab(!W_alu_result_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~2 .extended_lut = "off";
defparam \Equal1~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!W_alu_result_12),
	.datab(!W_alu_result_11),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~1 (
	.dataa(!W_alu_result_9),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal2),
	.datae(!\Equal4~0_combout ),
	.dataf(!\Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \Equal5~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~3 (
	.dataa(!Equal1),
	.datab(!Equal11),
	.datac(!Equal12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~3 .extended_lut = "off";
defparam \Equal1~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal1~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!W_alu_result_6),
	.datab(!W_alu_result_7),
	.datac(!W_alu_result_8),
	.datad(!W_alu_result_12),
	.datae(!W_alu_result_11),
	.dataf(!W_alu_result_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!W_alu_result_3),
	.datab(!W_alu_result_4),
	.datac(!W_alu_result_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal5~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_router_001 (
	F_pc_17,
	F_pc_16,
	F_pc_18,
	F_pc_19,
	F_pc_20,
	F_pc_21,
	F_pc_22,
	F_pc_23,
	F_pc_24,
	F_pc_26,
	F_pc_15,
	F_pc_14,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_25,
	Equal1,
	Equal11,
	Equal12,
	Equal2,
	Equal21,
	Equal13)/* synthesis synthesis_greybox=1 */;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_18;
input 	F_pc_19;
input 	F_pc_20;
input 	F_pc_21;
input 	F_pc_22;
input 	F_pc_23;
input 	F_pc_24;
input 	F_pc_26;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_9;
input 	F_pc_11;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_10;
input 	F_pc_25;
output 	Equal1;
output 	Equal11;
output 	Equal12;
output 	Equal2;
output 	Equal21;
output 	Equal13;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!F_pc_25),
	.datab(!F_pc_17),
	.datac(!F_pc_16),
	.datad(!F_pc_18),
	.datae(!F_pc_19),
	.dataf(!F_pc_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!F_pc_21),
	.datab(!F_pc_22),
	.datac(!F_pc_23),
	.datad(!F_pc_24),
	.datae(!F_pc_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~2 (
	.dataa(!F_pc_15),
	.datab(!F_pc_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~2 .extended_lut = "off";
defparam \Equal1~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!F_pc_15),
	.datab(!F_pc_14),
	.datac(!F_pc_11),
	.datad(!F_pc_13),
	.datae(!F_pc_12),
	.dataf(!F_pc_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!F_pc_9),
	.datab(!Equal2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~3 (
	.dataa(!Equal1),
	.datab(!Equal11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~3 .extended_lut = "off";
defparam \Equal1~3 .lut_mask = 64'h7777777777777777;
defparam \Equal1~3 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src1_valid,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src1_valid;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001_1 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_rsp_demux_001_2 (
	za_valid,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	za_valid;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!za_valid),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!za_valid),
	.datab(!mem_86_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_rsp_mux (
	ram_block1a32,
	ram_block1a0,
	av_readdata_pre_0,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a37,
	ram_block1a5,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	mem_86_0,
	mem_68_0,
	WideOr11,
	WideOr12,
	src0_valid2,
	av_readdata_pre_01,
	za_data_0,
	av_readdata_pre_02,
	address_reg_a_0,
	av_readdata_pre_03,
	src_data_0,
	za_data_24,
	av_readdata_pre_24,
	za_data_25,
	av_readdata_pre_25,
	za_data_26,
	av_readdata_pre_26,
	za_data_1,
	av_readdata_pre_11,
	za_data_4,
	av_readdata_pre_41,
	za_data_3,
	av_readdata_pre_31,
	za_data_2,
	av_readdata_pre_21,
	za_data_5,
	av_readdata_pre_51,
	za_data_28,
	av_readdata_pre_28,
	za_data_29,
	av_readdata_pre_29,
	za_data_30,
	av_readdata_pre_30,
	za_data_31,
	av_readdata_pre_311,
	za_data_27,
	av_readdata_pre_27,
	za_data_7,
	av_readdata_pre_71,
	za_data_6,
	av_readdata_pre_61,
	av_readdata_pre_12,
	av_readdata_pre_13,
	src_data_1,
	av_readdata_pre_22,
	av_readdata_pre_23,
	src_data_2,
	av_readdata_pre_32,
	av_readdata_pre_33,
	src_data_3,
	av_readdata_pre_42,
	av_readdata_pre_43,
	src_data_4,
	av_readdata_pre_52,
	av_readdata_pre_53,
	src_data_5,
	av_readdata_pre_62,
	av_readdata_pre_63,
	src_data_6,
	av_readdata_pre_72,
	av_readdata_pre_73,
	src_data_7,
	src_data_24,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31)/* synthesis synthesis_greybox=1 */;
input 	ram_block1a32;
input 	ram_block1a0;
input 	av_readdata_pre_0;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a38;
input 	ram_block1a6;
input 	av_readdata_pre_1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	mem_86_0;
input 	mem_68_0;
output 	WideOr11;
output 	WideOr12;
input 	src0_valid2;
input 	av_readdata_pre_01;
input 	za_data_0;
input 	av_readdata_pre_02;
input 	address_reg_a_0;
input 	av_readdata_pre_03;
output 	src_data_0;
input 	za_data_24;
input 	av_readdata_pre_24;
input 	za_data_25;
input 	av_readdata_pre_25;
input 	za_data_26;
input 	av_readdata_pre_26;
input 	za_data_1;
input 	av_readdata_pre_11;
input 	za_data_4;
input 	av_readdata_pre_41;
input 	za_data_3;
input 	av_readdata_pre_31;
input 	za_data_2;
input 	av_readdata_pre_21;
input 	za_data_5;
input 	av_readdata_pre_51;
input 	za_data_28;
input 	av_readdata_pre_28;
input 	za_data_29;
input 	av_readdata_pre_29;
input 	za_data_30;
input 	av_readdata_pre_30;
input 	za_data_31;
input 	av_readdata_pre_311;
input 	za_data_27;
input 	av_readdata_pre_27;
input 	za_data_7;
input 	av_readdata_pre_71;
input 	za_data_6;
input 	av_readdata_pre_61;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
output 	src_data_1;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
output 	src_data_2;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
output 	src_data_3;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
output 	src_data_4;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
output 	src_data_5;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
output 	src_data_6;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
output 	src_data_7;
output 	src_data_24;
output 	src_data_25;
output 	src_data_26;
output 	src_data_27;
output 	src_data_28;
output 	src_data_29;
output 	src_data_30;
output 	src_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_data[0]~24_combout ;
wire \src_data[0]~0_combout ;
wire \src_data[1]~25_combout ;
wire \src_data[1]~2_combout ;
wire \src_data[2]~26_combout ;
wire \src_data[2]~4_combout ;
wire \src_data[3]~27_combout ;
wire \src_data[3]~6_combout ;
wire \src_data[4]~28_combout ;
wire \src_data[4]~8_combout ;
wire \src_data[5]~29_combout ;
wire \src_data[5]~10_combout ;
wire \src_data[6]~30_combout ;
wire \src_data[6]~12_combout ;
wire \src_data[7]~31_combout ;
wire \src_data[7]~14_combout ;
wire \src_data[24]~32_combout ;
wire \src_data[25]~33_combout ;
wire \src_data[26]~34_combout ;
wire \src_data[27]~35_combout ;
wire \src_data[28]~36_combout ;
wire \src_data[29]~37_combout ;
wire \src_data[30]~38_combout ;
wire \src_data[31]~39_combout ;


cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!read_latency_shift_reg_02),
	.datad(!read_latency_shift_reg_03),
	.datae(!mem_86_0),
	.dataf(!mem_68_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!WideOr11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr12),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_01),
	.datad(!za_data_0),
	.datae(!\src_data[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~3 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_11),
	.datad(!za_data_1),
	.datae(!\src_data[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~3 .extended_lut = "off";
defparam \src_data[1]~3 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~5 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_21),
	.datad(!za_data_2),
	.datae(!\src_data[2]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~5 .extended_lut = "off";
defparam \src_data[2]~5 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~7 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!za_data_3),
	.datae(!\src_data[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~7 .extended_lut = "off";
defparam \src_data[3]~7 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~9 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_41),
	.datad(!za_data_4),
	.datae(!\src_data[4]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~9 .extended_lut = "off";
defparam \src_data[4]~9 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[4]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~11 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_51),
	.datad(!za_data_5),
	.datae(!\src_data[5]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~11 .extended_lut = "off";
defparam \src_data[5]~11 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[5]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~13 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_61),
	.datad(!za_data_6),
	.datae(!\src_data[6]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~13 .extended_lut = "off";
defparam \src_data[6]~13 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[6]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~15 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_71),
	.datad(!za_data_7),
	.datae(!\src_data[7]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~15 .extended_lut = "off";
defparam \src_data[7]~15 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[7]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~16 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a56),
	.datad(!ram_block1a24),
	.datae(!\src_data[24]~32_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~16 .extended_lut = "off";
defparam \src_data[24]~16 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[24]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~17 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a57),
	.datad(!ram_block1a25),
	.datae(!\src_data[25]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~17 .extended_lut = "off";
defparam \src_data[25]~17 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[25]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~18 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a58),
	.datad(!ram_block1a26),
	.datae(!\src_data[26]~34_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~18 .extended_lut = "off";
defparam \src_data[26]~18 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[26]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~19 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a59),
	.datad(!ram_block1a27),
	.datae(!\src_data[27]~35_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~19 .extended_lut = "off";
defparam \src_data[27]~19 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[27]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~20 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a60),
	.datad(!ram_block1a28),
	.datae(!\src_data[28]~36_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~20 .extended_lut = "off";
defparam \src_data[28]~20 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[28]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~21 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a61),
	.datad(!ram_block1a29),
	.datae(!\src_data[29]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~21 .extended_lut = "off";
defparam \src_data[29]~21 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[29]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~22 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a62),
	.datad(!ram_block1a30),
	.datae(!\src_data[30]~38_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~22 .extended_lut = "off";
defparam \src_data[30]~22 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[30]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~23 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a63),
	.datad(!ram_block1a31),
	.datae(!\src_data[31]~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~23 .extended_lut = "off";
defparam \src_data[31]~23 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \src_data[31]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~24 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_02),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_0),
	.dataf(!av_readdata_pre_03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~24 .extended_lut = "off";
defparam \src_data[0]~24 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[0]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!src0_valid),
	.datab(!ram_block1a32),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a0),
	.datae(!\src_data[0]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'hFFACFFFFFFACFFFF;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~25 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_12),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_1),
	.dataf(!av_readdata_pre_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~25 .extended_lut = "off";
defparam \src_data[1]~25 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[1]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~2 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a33),
	.datad(!ram_block1a1),
	.datae(!\src_data[1]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~2 .extended_lut = "off";
defparam \src_data[1]~2 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~26 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_22),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_2),
	.dataf(!av_readdata_pre_23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~26 .extended_lut = "off";
defparam \src_data[2]~26 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[2]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~4 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a34),
	.datad(!ram_block1a2),
	.datae(!\src_data[2]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~4 .extended_lut = "off";
defparam \src_data[2]~4 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~27 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_32),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_3),
	.dataf(!av_readdata_pre_33),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~27 .extended_lut = "off";
defparam \src_data[3]~27 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[3]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~6 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a35),
	.datad(!ram_block1a3),
	.datae(!\src_data[3]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~6 .extended_lut = "off";
defparam \src_data[3]~6 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~28 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_42),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_4),
	.dataf(!av_readdata_pre_43),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~28 .extended_lut = "off";
defparam \src_data[4]~28 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[4]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~8 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a36),
	.datad(!ram_block1a4),
	.datae(!\src_data[4]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~8 .extended_lut = "off";
defparam \src_data[4]~8 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~29 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_52),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_5),
	.dataf(!av_readdata_pre_53),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~29 .extended_lut = "off";
defparam \src_data[5]~29 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[5]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~10 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a37),
	.datad(!ram_block1a5),
	.datae(!\src_data[5]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~10 .extended_lut = "off";
defparam \src_data[5]~10 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~30 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_62),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_6),
	.dataf(!av_readdata_pre_63),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~30 .extended_lut = "off";
defparam \src_data[6]~30 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[6]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~12 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a38),
	.datad(!ram_block1a6),
	.datae(!\src_data[6]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~12 .extended_lut = "off";
defparam \src_data[6]~12 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[6]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~31 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_72),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg_01),
	.datae(!av_readdata_pre_7),
	.dataf(!av_readdata_pre_73),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~31 .extended_lut = "off";
defparam \src_data[7]~31 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \src_data[7]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~14 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a39),
	.datad(!ram_block1a7),
	.datae(!\src_data[7]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~14 .extended_lut = "off";
defparam \src_data[7]~14 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \src_data[7]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~32 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!za_data_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~32 .extended_lut = "off";
defparam \src_data[24]~32 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~33 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_25),
	.datad(!za_data_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~33 .extended_lut = "off";
defparam \src_data[25]~33 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[25]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~34 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!za_data_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~34 .extended_lut = "off";
defparam \src_data[26]~34 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[26]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~35 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_27),
	.datad(!za_data_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~35 .extended_lut = "off";
defparam \src_data[27]~35 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[27]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~36 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_28),
	.datad(!za_data_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~36 .extended_lut = "off";
defparam \src_data[28]~36 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[28]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~37 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!za_data_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[29]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~37 .extended_lut = "off";
defparam \src_data[29]~37 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~38 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_30),
	.datad(!za_data_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~38 .extended_lut = "off";
defparam \src_data[30]~38 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[30]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~39 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_311),
	.datad(!za_data_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~39 .extended_lut = "off";
defparam \src_data[31]~39 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[31]~39 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_mm_interconnect_0_rsp_mux_001 (
	src1_valid,
	src1_valid1,
	src1_valid2,
	WideOr1)/* synthesis synthesis_greybox=1 */;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
output 	WideOr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr1),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \WideOr1~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_24,
	W_alu_result_25,
	W_alu_result_26,
	W_alu_result_27,
	W_alu_result_28,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_21,
	W_alu_result_22,
	W_alu_result_23,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_17,
	F_pc_16,
	F_pc_18,
	F_pc_19,
	F_pc_20,
	F_pc_21,
	F_pc_22,
	F_pc_23,
	F_pc_24,
	F_pc_26,
	F_pc_15,
	F_pc_14,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	ram_block1a32,
	ram_block1a0,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a37,
	ram_block1a5,
	ram_block1a40,
	ram_block1a8,
	ram_block1a42,
	ram_block1a10,
	ram_block1a41,
	ram_block1a9,
	ram_block1a60,
	ram_block1a28,
	ram_block1a53,
	ram_block1a21,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	ram_block1a52,
	ram_block1a20,
	ram_block1a51,
	ram_block1a19,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	readdata_0,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_5,
	readdata_8,
	readdata_10,
	readdata_9,
	readdata_28,
	readdata_21,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_17,
	readdata_18,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_21,
	av_readdata_pre_22,
	readdata_27,
	av_readdata_pre_18,
	av_readdata_pre_17,
	readdata_7,
	readdata_6,
	av_readdata_pre_16,
	readdata_20,
	readdata_19,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write,
	always0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_read,
	av_waitrequest,
	sink_ready,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	WideOr0,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	av_waitrequest1,
	i_read,
	F_pc_25,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	rf_source_valid,
	src1_valid,
	src1_valid1,
	src1_valid2,
	WideOr12,
	hbreak_enabled,
	src0_valid2,
	av_readdata_pre_0,
	za_data_0,
	address_reg_a_0,
	src_data_0,
	za_data_22,
	av_readdata_pre_221,
	za_data_23,
	av_readdata_pre_23,
	za_data_24,
	av_readdata_pre_24,
	za_data_25,
	av_readdata_pre_25,
	za_data_26,
	av_readdata_pre_26,
	za_data_1,
	av_readdata_pre_1,
	za_data_4,
	av_readdata_pre_4,
	za_data_3,
	av_readdata_pre_3,
	za_data_2,
	av_readdata_pre_2,
	WideOr13,
	src_data_46,
	av_readdata_pre_11,
	za_data_11,
	za_data_12,
	av_readdata_pre_12,
	za_data_13,
	av_readdata_pre_13,
	za_data_14,
	av_readdata_pre_14,
	za_data_15,
	av_readdata_pre_15,
	za_data_16,
	av_readdata_pre_161,
	za_data_5,
	av_readdata_pre_5,
	za_data_8,
	av_readdata_pre_8,
	za_data_10,
	av_readdata_pre_10,
	za_data_9,
	av_readdata_pre_9,
	za_data_28,
	av_readdata_pre_28,
	za_data_21,
	av_readdata_pre_211,
	za_data_29,
	av_readdata_pre_29,
	za_data_30,
	av_readdata_pre_30,
	za_data_31,
	av_readdata_pre_31,
	za_data_17,
	av_readdata_pre_171,
	za_data_18,
	av_readdata_pre_181,
	za_data_27,
	av_readdata_pre_27,
	za_data_7,
	av_readdata_pre_7,
	za_data_6,
	av_readdata_pre_6,
	za_data_20,
	av_readdata_pre_201,
	za_data_19,
	av_readdata_pre_191,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	r_early_rst,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	av_readdata_pre_81,
	av_readdata_9,
	av_readdata_8,
	av_readdata_pre_91,
	src_data_24,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	av_readdata_pre_151,
	av_readdata_pre_141,
	av_readdata_pre_131,
	av_readdata_pre_121,
	av_readdata_pre_101,
	src_payload,
	src_data_38,
	src_data_40,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_41,
	src_payload1,
	src_data_32,
	src_data_29,
	src_data_30,
	src_data_31,
	src_payload2,
	src_payload3,
	debug_reset_request,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_33,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_9;
output 	W_alu_result_24;
output 	W_alu_result_25;
output 	W_alu_result_26;
output 	W_alu_result_27;
output 	W_alu_result_28;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_21;
output 	W_alu_result_22;
output 	W_alu_result_23;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_6;
output 	W_alu_result_7;
output 	W_alu_result_8;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_2;
output 	W_alu_result_3;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_18;
output 	F_pc_19;
output 	F_pc_20;
output 	F_pc_21;
output 	F_pc_22;
output 	F_pc_23;
output 	F_pc_24;
output 	F_pc_26;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_9;
output 	F_pc_11;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_10;
output 	F_pc_0;
output 	F_pc_1;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_7;
output 	F_pc_8;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a54;
input 	ram_block1a22;
input 	ram_block1a55;
input 	ram_block1a23;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a48;
input 	ram_block1a16;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a53;
input 	ram_block1a21;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	ram_block1a49;
input 	ram_block1a17;
input 	ram_block1a50;
input 	ram_block1a18;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a38;
input 	ram_block1a6;
input 	ram_block1a52;
input 	ram_block1a20;
input 	ram_block1a51;
input 	ram_block1a19;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
output 	readdata_0;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_5;
output 	readdata_8;
output 	readdata_10;
output 	readdata_9;
output 	readdata_28;
output 	readdata_21;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
output 	readdata_17;
output 	readdata_18;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
output 	readdata_27;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
output 	readdata_7;
output 	readdata_6;
input 	av_readdata_pre_16;
output 	readdata_20;
output 	readdata_19;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write;
input 	always0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_read;
input 	av_waitrequest;
input 	sink_ready;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	WideOr0;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	WideOr11;
input 	av_waitrequest1;
output 	i_read;
output 	F_pc_25;
output 	d_byteenable_0;
output 	d_byteenable_1;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	rf_source_valid;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	WideOr12;
output 	hbreak_enabled;
input 	src0_valid2;
input 	av_readdata_pre_0;
input 	za_data_0;
input 	address_reg_a_0;
input 	src_data_0;
input 	za_data_22;
input 	av_readdata_pre_221;
input 	za_data_23;
input 	av_readdata_pre_23;
input 	za_data_24;
input 	av_readdata_pre_24;
input 	za_data_25;
input 	av_readdata_pre_25;
input 	za_data_26;
input 	av_readdata_pre_26;
input 	za_data_1;
input 	av_readdata_pre_1;
input 	za_data_4;
input 	av_readdata_pre_4;
input 	za_data_3;
input 	av_readdata_pre_3;
input 	za_data_2;
input 	av_readdata_pre_2;
input 	WideOr13;
input 	src_data_46;
input 	av_readdata_pre_11;
input 	za_data_11;
input 	za_data_12;
input 	av_readdata_pre_12;
input 	za_data_13;
input 	av_readdata_pre_13;
input 	za_data_14;
input 	av_readdata_pre_14;
input 	za_data_15;
input 	av_readdata_pre_15;
input 	za_data_16;
input 	av_readdata_pre_161;
input 	za_data_5;
input 	av_readdata_pre_5;
input 	za_data_8;
input 	av_readdata_pre_8;
input 	za_data_10;
input 	av_readdata_pre_10;
input 	za_data_9;
input 	av_readdata_pre_9;
input 	za_data_28;
input 	av_readdata_pre_28;
input 	za_data_21;
input 	av_readdata_pre_211;
input 	za_data_29;
input 	av_readdata_pre_29;
input 	za_data_30;
input 	av_readdata_pre_30;
input 	za_data_31;
input 	av_readdata_pre_31;
input 	za_data_17;
input 	av_readdata_pre_171;
input 	za_data_18;
input 	av_readdata_pre_181;
input 	za_data_27;
input 	av_readdata_pre_27;
input 	za_data_7;
input 	av_readdata_pre_7;
input 	za_data_6;
input 	av_readdata_pre_6;
input 	za_data_20;
input 	av_readdata_pre_201;
input 	za_data_19;
input 	av_readdata_pre_191;
input 	src_data_1;
input 	src_data_2;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	r_early_rst;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	av_readdata_pre_81;
input 	av_readdata_9;
input 	av_readdata_8;
input 	av_readdata_pre_91;
input 	src_data_24;
input 	src_data_25;
input 	src_data_26;
input 	src_data_27;
input 	src_data_28;
input 	av_readdata_pre_151;
input 	av_readdata_pre_141;
input 	av_readdata_pre_131;
input 	av_readdata_pre_121;
input 	av_readdata_pre_101;
input 	src_payload;
input 	src_data_38;
input 	src_data_40;
input 	src_data_39;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_data_41;
input 	src_payload1;
input 	src_data_32;
input 	src_data_29;
input 	src_data_30;
input 	src_data_31;
input 	src_payload2;
input 	src_payload3;
output 	debug_reset_request;
input 	src_payload4;
input 	src_payload5;
input 	src_data_34;
input 	src_payload6;
input 	src_payload7;
input 	src_data_35;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_data_33;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_sdram_demo_nios2_cpu cpu(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_18(F_pc_18),
	.F_pc_19(F_pc_19),
	.F_pc_20(F_pc_20),
	.F_pc_21(F_pc_21),
	.F_pc_22(F_pc_22),
	.F_pc_23(F_pc_23),
	.F_pc_24(F_pc_24),
	.F_pc_26(F_pc_26),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_9(F_pc_9),
	.F_pc_11(F_pc_11),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_10(F_pc_10),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.F_pc_8(F_pc_8),
	.ram_block1a32(ram_block1a32),
	.ram_block1a0(ram_block1a0),
	.ram_block1a54(ram_block1a54),
	.ram_block1a22(ram_block1a22),
	.ram_block1a55(ram_block1a55),
	.ram_block1a23(ram_block1a23),
	.ram_block1a56(ram_block1a56),
	.ram_block1a24(ram_block1a24),
	.ram_block1a57(ram_block1a57),
	.ram_block1a25(ram_block1a25),
	.ram_block1a58(ram_block1a58),
	.ram_block1a26(ram_block1a26),
	.ram_block1a33(ram_block1a33),
	.ram_block1a1(ram_block1a1),
	.ram_block1a36(ram_block1a36),
	.ram_block1a4(ram_block1a4),
	.ram_block1a35(ram_block1a35),
	.ram_block1a3(ram_block1a3),
	.ram_block1a34(ram_block1a34),
	.ram_block1a2(ram_block1a2),
	.ram_block1a43(ram_block1a43),
	.ram_block1a11(ram_block1a11),
	.ram_block1a44(ram_block1a44),
	.ram_block1a12(ram_block1a12),
	.ram_block1a45(ram_block1a45),
	.ram_block1a13(ram_block1a13),
	.ram_block1a46(ram_block1a46),
	.ram_block1a14(ram_block1a14),
	.ram_block1a47(ram_block1a47),
	.ram_block1a15(ram_block1a15),
	.ram_block1a48(ram_block1a48),
	.ram_block1a16(ram_block1a16),
	.ram_block1a37(ram_block1a37),
	.ram_block1a5(ram_block1a5),
	.ram_block1a40(ram_block1a40),
	.ram_block1a8(ram_block1a8),
	.ram_block1a42(ram_block1a42),
	.ram_block1a10(ram_block1a10),
	.ram_block1a41(ram_block1a41),
	.ram_block1a9(ram_block1a9),
	.ram_block1a60(ram_block1a60),
	.ram_block1a28(ram_block1a28),
	.ram_block1a53(ram_block1a53),
	.ram_block1a21(ram_block1a21),
	.ram_block1a61(ram_block1a61),
	.ram_block1a29(ram_block1a29),
	.ram_block1a62(ram_block1a62),
	.ram_block1a30(ram_block1a30),
	.ram_block1a63(ram_block1a63),
	.ram_block1a31(ram_block1a31),
	.ram_block1a49(ram_block1a49),
	.ram_block1a17(ram_block1a17),
	.ram_block1a50(ram_block1a50),
	.ram_block1a18(ram_block1a18),
	.ram_block1a59(ram_block1a59),
	.ram_block1a27(ram_block1a27),
	.ram_block1a39(ram_block1a39),
	.ram_block1a7(ram_block1a7),
	.ram_block1a38(ram_block1a38),
	.ram_block1a6(ram_block1a6),
	.ram_block1a52(ram_block1a52),
	.ram_block1a20(ram_block1a20),
	.ram_block1a51(ram_block1a51),
	.ram_block1a19(ram_block1a19),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.readdata_0(readdata_0),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_1(readdata_1),
	.readdata_4(readdata_4),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.readdata_11(readdata_11),
	.readdata_12(readdata_12),
	.readdata_13(readdata_13),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_16(readdata_16),
	.readdata_5(readdata_5),
	.readdata_8(readdata_8),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_28(readdata_28),
	.readdata_21(readdata_21),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.readdata_17(readdata_17),
	.readdata_18(readdata_18),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.readdata_27(readdata_27),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.av_readdata_pre_16(av_readdata_pre_16),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_write1(d_write),
	.always0(always0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_read1(d_read),
	.av_waitrequest(av_waitrequest),
	.sink_ready(sink_ready),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr0(WideOr0),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.WideOr1(WideOr1),
	.WideOr11(WideOr11),
	.av_waitrequest1(av_waitrequest1),
	.i_read1(i_read),
	.F_pc_25(F_pc_25),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.rf_source_valid(rf_source_valid),
	.src1_valid(src1_valid),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.WideOr12(WideOr12),
	.hbreak_enabled1(hbreak_enabled),
	.src0_valid2(src0_valid2),
	.av_readdata_pre_0(av_readdata_pre_0),
	.za_data_0(za_data_0),
	.address_reg_a_0(address_reg_a_0),
	.src_data_0(src_data_0),
	.za_data_22(za_data_22),
	.av_readdata_pre_221(av_readdata_pre_221),
	.za_data_23(za_data_23),
	.av_readdata_pre_23(av_readdata_pre_23),
	.za_data_24(za_data_24),
	.av_readdata_pre_24(av_readdata_pre_24),
	.za_data_25(za_data_25),
	.av_readdata_pre_25(av_readdata_pre_25),
	.za_data_26(za_data_26),
	.av_readdata_pre_26(av_readdata_pre_26),
	.za_data_1(za_data_1),
	.av_readdata_pre_1(av_readdata_pre_1),
	.za_data_4(za_data_4),
	.av_readdata_pre_4(av_readdata_pre_4),
	.za_data_3(za_data_3),
	.av_readdata_pre_3(av_readdata_pre_3),
	.za_data_2(za_data_2),
	.av_readdata_pre_2(av_readdata_pre_2),
	.WideOr13(WideOr13),
	.src_data_46(src_data_46),
	.av_readdata_pre_11(av_readdata_pre_11),
	.za_data_11(za_data_11),
	.za_data_12(za_data_12),
	.av_readdata_pre_12(av_readdata_pre_12),
	.za_data_13(za_data_13),
	.av_readdata_pre_13(av_readdata_pre_13),
	.za_data_14(za_data_14),
	.av_readdata_pre_14(av_readdata_pre_14),
	.za_data_15(za_data_15),
	.av_readdata_pre_15(av_readdata_pre_15),
	.za_data_16(za_data_16),
	.av_readdata_pre_161(av_readdata_pre_161),
	.za_data_5(za_data_5),
	.av_readdata_pre_5(av_readdata_pre_5),
	.za_data_8(za_data_8),
	.av_readdata_pre_8(av_readdata_pre_8),
	.za_data_10(za_data_10),
	.av_readdata_pre_10(av_readdata_pre_10),
	.za_data_9(za_data_9),
	.av_readdata_pre_9(av_readdata_pre_9),
	.za_data_28(za_data_28),
	.av_readdata_pre_28(av_readdata_pre_28),
	.za_data_21(za_data_21),
	.av_readdata_pre_211(av_readdata_pre_211),
	.za_data_29(za_data_29),
	.av_readdata_pre_29(av_readdata_pre_29),
	.za_data_30(za_data_30),
	.av_readdata_pre_30(av_readdata_pre_30),
	.za_data_31(za_data_31),
	.av_readdata_pre_31(av_readdata_pre_31),
	.za_data_17(za_data_17),
	.av_readdata_pre_171(av_readdata_pre_171),
	.za_data_18(za_data_18),
	.av_readdata_pre_181(av_readdata_pre_181),
	.za_data_27(za_data_27),
	.av_readdata_pre_27(av_readdata_pre_27),
	.za_data_7(za_data_7),
	.av_readdata_pre_7(av_readdata_pre_7),
	.za_data_6(za_data_6),
	.av_readdata_pre_6(av_readdata_pre_6),
	.za_data_20(za_data_20),
	.av_readdata_pre_201(av_readdata_pre_201),
	.za_data_19(za_data_19),
	.av_readdata_pre_191(av_readdata_pre_191),
	.src_data_1(src_data_1),
	.src_data_2(src_data_2),
	.src_data_3(src_data_3),
	.src_data_4(src_data_4),
	.src_data_5(src_data_5),
	.src_data_6(src_data_6),
	.src_data_7(src_data_7),
	.r_early_rst(r_early_rst),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.av_readdata_pre_81(av_readdata_pre_81),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.av_readdata_pre_91(av_readdata_pre_91),
	.src_data_24(src_data_24),
	.src_data_25(src_data_25),
	.src_data_26(src_data_26),
	.src_data_27(src_data_27),
	.src_data_28(src_data_28),
	.av_readdata_pre_151(av_readdata_pre_151),
	.av_readdata_pre_141(av_readdata_pre_141),
	.av_readdata_pre_131(av_readdata_pre_131),
	.av_readdata_pre_121(av_readdata_pre_121),
	.av_readdata_pre_101(av_readdata_pre_101),
	.src_payload(src_payload),
	.src_data_38(src_data_38),
	.src_data_40(src_data_40),
	.src_data_39(src_data_39),
	.src_data_45(src_data_45),
	.src_data_44(src_data_44),
	.src_data_43(src_data_43),
	.src_data_42(src_data_42),
	.src_data_41(src_data_41),
	.src_payload1(src_payload1),
	.src_data_32(src_data_32),
	.src_data_29(src_data_29),
	.src_data_30(src_data_30),
	.src_data_31(src_data_31),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.debug_reset_request(debug_reset_request),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_data_34(src_data_34),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_data_35(src_data_35),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_data_33(src_data_33),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module sdram_demo_sdram_demo_nios2_cpu (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_9,
	W_alu_result_24,
	W_alu_result_25,
	W_alu_result_26,
	W_alu_result_27,
	W_alu_result_28,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_21,
	W_alu_result_22,
	W_alu_result_23,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_8,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_2,
	W_alu_result_3,
	F_pc_17,
	F_pc_16,
	F_pc_18,
	F_pc_19,
	F_pc_20,
	F_pc_21,
	F_pc_22,
	F_pc_23,
	F_pc_24,
	F_pc_26,
	F_pc_15,
	F_pc_14,
	F_pc_9,
	F_pc_11,
	F_pc_13,
	F_pc_12,
	F_pc_10,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	F_pc_8,
	ram_block1a32,
	ram_block1a0,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a37,
	ram_block1a5,
	ram_block1a40,
	ram_block1a8,
	ram_block1a42,
	ram_block1a10,
	ram_block1a41,
	ram_block1a9,
	ram_block1a60,
	ram_block1a28,
	ram_block1a53,
	ram_block1a21,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	ram_block1a52,
	ram_block1a20,
	ram_block1a51,
	ram_block1a19,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	readdata_0,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_5,
	readdata_8,
	readdata_10,
	readdata_9,
	readdata_28,
	readdata_21,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_17,
	readdata_18,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_21,
	av_readdata_pre_22,
	readdata_27,
	av_readdata_pre_18,
	av_readdata_pre_17,
	readdata_7,
	readdata_6,
	av_readdata_pre_16,
	readdata_20,
	readdata_19,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write1,
	always0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_read1,
	av_waitrequest,
	sink_ready,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	WideOr0,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_0,
	WideOr1,
	WideOr11,
	av_waitrequest1,
	i_read1,
	F_pc_25,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	rf_source_valid,
	src1_valid,
	src1_valid1,
	src1_valid2,
	WideOr12,
	hbreak_enabled1,
	src0_valid2,
	av_readdata_pre_0,
	za_data_0,
	address_reg_a_0,
	src_data_0,
	za_data_22,
	av_readdata_pre_221,
	za_data_23,
	av_readdata_pre_23,
	za_data_24,
	av_readdata_pre_24,
	za_data_25,
	av_readdata_pre_25,
	za_data_26,
	av_readdata_pre_26,
	za_data_1,
	av_readdata_pre_1,
	za_data_4,
	av_readdata_pre_4,
	za_data_3,
	av_readdata_pre_3,
	za_data_2,
	av_readdata_pre_2,
	WideOr13,
	src_data_46,
	av_readdata_pre_11,
	za_data_11,
	za_data_12,
	av_readdata_pre_12,
	za_data_13,
	av_readdata_pre_13,
	za_data_14,
	av_readdata_pre_14,
	za_data_15,
	av_readdata_pre_15,
	za_data_16,
	av_readdata_pre_161,
	za_data_5,
	av_readdata_pre_5,
	za_data_8,
	av_readdata_pre_8,
	za_data_10,
	av_readdata_pre_10,
	za_data_9,
	av_readdata_pre_9,
	za_data_28,
	av_readdata_pre_28,
	za_data_21,
	av_readdata_pre_211,
	za_data_29,
	av_readdata_pre_29,
	za_data_30,
	av_readdata_pre_30,
	za_data_31,
	av_readdata_pre_31,
	za_data_17,
	av_readdata_pre_171,
	za_data_18,
	av_readdata_pre_181,
	za_data_27,
	av_readdata_pre_27,
	za_data_7,
	av_readdata_pre_7,
	za_data_6,
	av_readdata_pre_6,
	za_data_20,
	av_readdata_pre_201,
	za_data_19,
	av_readdata_pre_191,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	r_early_rst,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	av_readdata_pre_81,
	av_readdata_9,
	av_readdata_8,
	av_readdata_pre_91,
	src_data_24,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	av_readdata_pre_151,
	av_readdata_pre_141,
	av_readdata_pre_131,
	av_readdata_pre_121,
	av_readdata_pre_101,
	src_payload,
	src_data_38,
	src_data_40,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_41,
	src_payload1,
	src_data_32,
	src_data_29,
	src_data_30,
	src_data_31,
	src_payload2,
	src_payload3,
	debug_reset_request,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_33,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_9;
output 	W_alu_result_24;
output 	W_alu_result_25;
output 	W_alu_result_26;
output 	W_alu_result_27;
output 	W_alu_result_28;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_21;
output 	W_alu_result_22;
output 	W_alu_result_23;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_6;
output 	W_alu_result_7;
output 	W_alu_result_8;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_2;
output 	W_alu_result_3;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_18;
output 	F_pc_19;
output 	F_pc_20;
output 	F_pc_21;
output 	F_pc_22;
output 	F_pc_23;
output 	F_pc_24;
output 	F_pc_26;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_9;
output 	F_pc_11;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_10;
output 	F_pc_0;
output 	F_pc_1;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_7;
output 	F_pc_8;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a54;
input 	ram_block1a22;
input 	ram_block1a55;
input 	ram_block1a23;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a48;
input 	ram_block1a16;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a53;
input 	ram_block1a21;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	ram_block1a49;
input 	ram_block1a17;
input 	ram_block1a50;
input 	ram_block1a18;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a38;
input 	ram_block1a6;
input 	ram_block1a52;
input 	ram_block1a20;
input 	ram_block1a51;
input 	ram_block1a19;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
output 	readdata_0;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_5;
output 	readdata_8;
output 	readdata_10;
output 	readdata_9;
output 	readdata_28;
output 	readdata_21;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
output 	readdata_17;
output 	readdata_18;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
output 	readdata_27;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
output 	readdata_7;
output 	readdata_6;
input 	av_readdata_pre_16;
output 	readdata_20;
output 	readdata_19;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write1;
input 	always0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_read1;
input 	av_waitrequest;
input 	sink_ready;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	WideOr0;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	WideOr11;
input 	av_waitrequest1;
output 	i_read1;
output 	F_pc_25;
output 	d_byteenable_0;
output 	d_byteenable_1;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	rf_source_valid;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	WideOr12;
output 	hbreak_enabled1;
input 	src0_valid2;
input 	av_readdata_pre_0;
input 	za_data_0;
input 	address_reg_a_0;
input 	src_data_0;
input 	za_data_22;
input 	av_readdata_pre_221;
input 	za_data_23;
input 	av_readdata_pre_23;
input 	za_data_24;
input 	av_readdata_pre_24;
input 	za_data_25;
input 	av_readdata_pre_25;
input 	za_data_26;
input 	av_readdata_pre_26;
input 	za_data_1;
input 	av_readdata_pre_1;
input 	za_data_4;
input 	av_readdata_pre_4;
input 	za_data_3;
input 	av_readdata_pre_3;
input 	za_data_2;
input 	av_readdata_pre_2;
input 	WideOr13;
input 	src_data_46;
input 	av_readdata_pre_11;
input 	za_data_11;
input 	za_data_12;
input 	av_readdata_pre_12;
input 	za_data_13;
input 	av_readdata_pre_13;
input 	za_data_14;
input 	av_readdata_pre_14;
input 	za_data_15;
input 	av_readdata_pre_15;
input 	za_data_16;
input 	av_readdata_pre_161;
input 	za_data_5;
input 	av_readdata_pre_5;
input 	za_data_8;
input 	av_readdata_pre_8;
input 	za_data_10;
input 	av_readdata_pre_10;
input 	za_data_9;
input 	av_readdata_pre_9;
input 	za_data_28;
input 	av_readdata_pre_28;
input 	za_data_21;
input 	av_readdata_pre_211;
input 	za_data_29;
input 	av_readdata_pre_29;
input 	za_data_30;
input 	av_readdata_pre_30;
input 	za_data_31;
input 	av_readdata_pre_31;
input 	za_data_17;
input 	av_readdata_pre_171;
input 	za_data_18;
input 	av_readdata_pre_181;
input 	za_data_27;
input 	av_readdata_pre_27;
input 	za_data_7;
input 	av_readdata_pre_7;
input 	za_data_6;
input 	av_readdata_pre_6;
input 	za_data_20;
input 	av_readdata_pre_201;
input 	za_data_19;
input 	av_readdata_pre_191;
input 	src_data_1;
input 	src_data_2;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	r_early_rst;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	av_readdata_pre_81;
input 	av_readdata_9;
input 	av_readdata_8;
input 	av_readdata_pre_91;
input 	src_data_24;
input 	src_data_25;
input 	src_data_26;
input 	src_data_27;
input 	src_data_28;
input 	av_readdata_pre_151;
input 	av_readdata_pre_141;
input 	av_readdata_pre_131;
input 	av_readdata_pre_121;
input 	av_readdata_pre_101;
input 	src_payload;
input 	src_data_38;
input 	src_data_40;
input 	src_data_39;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_data_41;
input 	src_payload1;
input 	src_data_32;
input 	src_data_29;
input 	src_data_30;
input 	src_data_31;
input 	src_payload2;
input 	src_payload3;
output 	debug_reset_request;
input 	src_payload4;
input 	src_payload5;
input 	src_data_34;
input 	src_payload6;
input 	src_payload7;
input 	src_data_35;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_data_33;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \av_ld_byte0_data[0]~q ;
wire \W_alu_result[0]~q ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \av_ld_byte0_data[1]~q ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte0_data[2]~q ;
wire \av_ld_byte0_data[3]~q ;
wire \av_ld_byte0_data[4]~q ;
wire \av_ld_byte0_data[5]~q ;
wire \av_ld_byte0_data[6]~q ;
wire \av_ld_byte0_data[7]~q ;
wire \av_ld_byte3_data[0]~q ;
wire \av_ld_byte3_data[1]~q ;
wire \av_ld_byte3_data[2]~q ;
wire \av_ld_byte3_data[3]~q ;
wire \av_ld_byte3_data[4]~q ;
wire \Add2~125_sumout ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \av_ld_byte3_data[5]~q ;
wire \av_ld_byte3_data[6]~q ;
wire \av_ld_byte3_data[7]~q ;
wire \Add2~129_sumout ;
wire \W_alu_result[31]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[29]~q ;
wire \Add2~133_sumout ;
wire \E_control_rd_data[0]~1_combout ;
wire \W_rf_wr_data[0]~31_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \W_control_rd_data[0]~q ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \W_rf_wr_data[1]~0_combout ;
wire \W_rf_wr_data[2]~1_combout ;
wire \W_rf_wr_data[3]~2_combout ;
wire \W_rf_wr_data[4]~3_combout ;
wire \W_rf_wr_data[5]~4_combout ;
wire \W_rf_wr_data[6]~5_combout ;
wire \W_rf_wr_data[7]~6_combout ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_dst_regnum[1]~1_combout ;
wire \D_dst_regnum[2]~2_combout ;
wire \D_dst_regnum[2]~3_combout ;
wire \D_dst_regnum[3]~4_combout ;
wire \D_dst_regnum[3]~5_combout ;
wire \D_dst_regnum[0]~6_combout ;
wire \D_dst_regnum[0]~7_combout ;
wire \D_dst_regnum[4]~8_combout ;
wire \D_dst_regnum[4]~9_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \D_ctrl_ld_signed~0_combout ;
wire \av_ld_byte1_data[0]~q ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_byte0_data[7]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_alu_result[0]~28_combout ;
wire \the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|jtag_break~q ;
wire \av_ld_byte1_data[1]~q ;
wire \W_rf_wr_data[9]~7_combout ;
wire \W_rf_wr_data[24]~8_combout ;
wire \W_rf_wr_data[25]~9_combout ;
wire \W_rf_wr_data[26]~10_combout ;
wire \W_rf_wr_data[27]~11_combout ;
wire \W_rf_wr_data[28]~12_combout ;
wire \av_ld_byte2_data[4]~q ;
wire \W_rf_wr_data[20]~13_combout ;
wire \av_ld_byte2_data[3]~q ;
wire \W_rf_wr_data[19]~14_combout ;
wire \av_ld_byte2_data[5]~q ;
wire \W_rf_wr_data[21]~15_combout ;
wire \av_ld_byte2_data[6]~q ;
wire \W_rf_wr_data[22]~16_combout ;
wire \av_ld_byte2_data[7]~q ;
wire \W_rf_wr_data[23]~17_combout ;
wire \av_ld_byte2_data[2]~q ;
wire \W_rf_wr_data[18]~18_combout ;
wire \av_ld_byte2_data[1]~q ;
wire \W_rf_wr_data[17]~19_combout ;
wire \av_ld_byte2_data[0]~q ;
wire \W_rf_wr_data[16]~20_combout ;
wire \av_ld_byte1_data[7]~q ;
wire \W_rf_wr_data[15]~21_combout ;
wire \av_ld_byte1_data[6]~q ;
wire \W_rf_wr_data[14]~22_combout ;
wire \av_ld_byte1_data[5]~q ;
wire \W_rf_wr_data[13]~23_combout ;
wire \W_rf_wr_data[8]~24_combout ;
wire \av_ld_byte1_data[4]~q ;
wire \W_rf_wr_data[12]~25_combout ;
wire \av_ld_byte1_data[3]~q ;
wire \W_rf_wr_data[11]~26_combout ;
wire \av_ld_byte1_data[2]~q ;
wire \W_rf_wr_data[10]~27_combout ;
wire \E_alu_result[1]~29_combout ;
wire \LessThan0~0_combout ;
wire \av_ld_byte1_data_nxt[0]~0_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_nxt[0]~1_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \av_ld_byte1_data_nxt[1]~2_combout ;
wire \av_ld_byte1_data_nxt[1]~3_combout ;
wire \av_ld_byte2_data_nxt[4]~0_combout ;
wire \av_ld_byte2_data_nxt[4]~1_combout ;
wire \av_ld_byte2_data_nxt[3]~2_combout ;
wire \av_ld_byte2_data_nxt[3]~3_combout ;
wire \av_ld_byte2_data_nxt[5]~4_combout ;
wire \av_ld_byte2_data_nxt[5]~5_combout ;
wire \av_ld_byte2_data_nxt[6]~6_combout ;
wire \av_ld_byte2_data_nxt[6]~7_combout ;
wire \av_ld_byte2_data_nxt[7]~8_combout ;
wire \av_ld_byte2_data_nxt[7]~9_combout ;
wire \av_ld_byte2_data_nxt[2]~10_combout ;
wire \av_ld_byte2_data_nxt[2]~11_combout ;
wire \av_ld_byte2_data_nxt[1]~12_combout ;
wire \av_ld_byte2_data_nxt[1]~13_combout ;
wire \av_ld_byte2_data_nxt[0]~14_combout ;
wire \av_ld_byte2_data_nxt[0]~15_combout ;
wire \av_ld_byte1_data_nxt[7]~4_combout ;
wire \av_ld_byte1_data_nxt[7]~5_combout ;
wire \av_ld_byte1_data_nxt[6]~6_combout ;
wire \av_ld_byte1_data_nxt[6]~7_combout ;
wire \av_ld_byte1_data_nxt[5]~8_combout ;
wire \av_ld_byte1_data_nxt[5]~9_combout ;
wire \av_ld_byte1_data_nxt[4]~10_combout ;
wire \av_ld_byte1_data_nxt[4]~11_combout ;
wire \av_ld_byte1_data_nxt[3]~12_combout ;
wire \av_ld_byte1_data_nxt[3]~13_combout ;
wire \av_ld_byte1_data_nxt[2]~14_combout ;
wire \av_ld_byte1_data_nxt[2]~15_combout ;
wire \W_rf_wr_data[31]~28_combout ;
wire \W_rf_wr_data[30]~29_combout ;
wire \W_rf_wr_data[29]~30_combout ;
wire \E_alu_result[31]~30_combout ;
wire \E_alu_result[30]~31_combout ;
wire \E_alu_result[29]~32_combout ;
wire \av_ld_byte1_data_nxt[0]~16_combout ;
wire \av_ld_byte1_data_nxt[4]~17_combout ;
wire \av_ld_byte1_data_nxt[3]~18_combout ;
wire \av_ld_byte1_data_nxt[2]~19_combout ;
wire \av_ld_byte1_data_nxt[1]~20_combout ;
wire \av_ld_byte2_data_nxt[1]~16_combout ;
wire \av_ld_byte2_data_nxt[0]~17_combout ;
wire \av_ld_byte1_data_nxt[7]~21_combout ;
wire \av_ld_byte1_data_nxt[6]~22_combout ;
wire \av_ld_byte1_data_nxt[5]~23_combout ;
wire \av_ld_byte2_data_nxt[4]~18_combout ;
wire \av_ld_byte2_data_nxt[3]~19_combout ;
wire \av_ld_byte2_data_nxt[5]~20_combout ;
wire \av_ld_byte2_data_nxt[6]~21_combout ;
wire \av_ld_byte2_data_nxt[7]~22_combout ;
wire \av_ld_byte2_data_nxt[2]~23_combout ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \F_iw[0]~41_combout ;
wire \F_iw[0]~5_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \E_new_inst~q ;
wire \F_iw[1]~57_combout ;
wire \F_iw[1]~6_combout ;
wire \D_iw[1]~q ;
wire \F_iw[4]~59_combout ;
wire \F_iw[4]~7_combout ;
wire \D_iw[4]~q ;
wire \F_iw[3]~58_combout ;
wire \F_iw[3]~8_combout ;
wire \D_iw[3]~q ;
wire \D_ctrl_st~0_combout ;
wire \F_iw[2]~42_combout ;
wire \F_iw[2]~9_combout ;
wire \D_iw[2]~q ;
wire \R_ctrl_st~q ;
wire \d_write_nxt~0_combout ;
wire \E_st_stall~combout ;
wire \D_ctrl_ld~0_combout ;
wire \R_ctrl_ld~q ;
wire \E_ld_stall~0_combout ;
wire \av_ld_aligning_data~q ;
wire \D_ctrl_mem16~0_combout ;
wire \av_ld_align_cycle_nxt[0]~1_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \av_ld_align_cycle_nxt[1]~0_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \E_stall~0_combout ;
wire \F_iw[6]~43_combout ;
wire \F_iw[6]~29_combout ;
wire \D_iw[6]~q ;
wire \F_iw[5]~60_combout ;
wire \F_iw[5]~16_combout ;
wire \D_iw[5]~q ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \F_iw[13]~54_combout ;
wire \F_iw[13]~12_combout ;
wire \D_iw[13]~q ;
wire \F_iw[12]~40_combout ;
wire \F_iw[12]~11_combout ;
wire \D_iw[12]~q ;
wire \F_iw[15]~55_combout ;
wire \F_iw[15]~14_combout ;
wire \D_iw[15]~q ;
wire \F_iw[11]~33_combout ;
wire \F_iw[11]~10_combout ;
wire \D_iw[11]~q ;
wire \F_iw[14]~34_combout ;
wire \F_iw[14]~13_combout ;
wire \D_iw[14]~q ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~5_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \R_src2_lo~0_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \Equal62~6_combout ;
wire \Equal62~7_combout ;
wire \D_ctrl_implicit_dst_eretaddr~6_combout ;
wire \D_ctrl_implicit_dst_eretaddr~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~4_combout ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \Equal0~12_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~8_combout ;
wire \Equal62~9_combout ;
wire \Equal62~10_combout ;
wire \Equal62~12_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal0~9_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \Equal0~13_combout ;
wire \Equal62~14_combout ;
wire \Equal62~15_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[0]~5_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~_wirecell_combout ;
wire \E_shift_rot_cnt[0]~q ;
wire \Add3~3_combout ;
wire \F_iw[7]~45_combout ;
wire \F_iw[7]~28_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~4_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \Add3~2_combout ;
wire \F_iw[8]~44_combout ;
wire \F_iw[8]~17_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~2_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \Add3~1_combout ;
wire \F_iw[9]~46_combout ;
wire \F_iw[9]~19_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~3_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_stall~1_combout ;
wire \Add3~0_combout ;
wire \F_iw[10]~47_combout ;
wire \F_iw[10]~18_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~1_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~2_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_valid_from_R~0_combout ;
wire \E_valid_from_R~q ;
wire \W_valid~0_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \D_iw[0]~q ;
wire \Equal0~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~3_combout ;
wire \Equal0~11_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~0_combout ;
wire \R_ctrl_exception~q ;
wire \D_ctrl_break~0_combout ;
wire \D_ctrl_break~1_combout ;
wire \R_ctrl_break~q ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~0_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_src1~1_combout ;
wire \R_src1[0]~33_combout ;
wire \E_src1[0]~q ;
wire \Equal132~1_combout ;
wire \Equal133~0_combout ;
wire \Equal62~16_combout ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \W_estatus_reg~q ;
wire \Equal134~0_combout ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \W_bstatus_reg~q ;
wire \Equal132~0_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \Equal135~0_combout ;
wire \W_ienable_reg[0]~0_combout ;
wire \W_ienable_reg[0]~q ;
wire \W_ipending_reg_nxt[0]~0_combout ;
wire \W_ipending_reg[0]~q ;
wire \intr_req~combout ;
wire \D_iw[1]~0_combout ;
wire \F_iw[16]~56_combout ;
wire \F_iw[16]~15_combout ;
wire \D_iw[16]~q ;
wire \D_ctrl_shift_rot~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \R_ctrl_shift_rot~q ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~1_combout ;
wire \R_ctrl_logic~q ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \Equal62~0_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \R_ctrl_shift_logical~q ;
wire \Equal62~1_combout ;
wire \R_ctrl_rot_right_nxt~combout ;
wire \R_ctrl_rot_right~q ;
wire \E_shift_rot_result_nxt[5]~1_combout ;
wire \Add0~102 ;
wire \Add0~106 ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \R_src1[5]~3_combout ;
wire \E_src1[5]~q ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[6]~19_combout ;
wire \Add0~6 ;
wire \Add0~77_sumout ;
wire \R_src1[6]~21_combout ;
wire \E_src1[6]~q ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[7]~20_combout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \R_src1[7]~22_combout ;
wire \E_src1[7]~q ;
wire \E_shift_rot_result[7]~q ;
wire \E_shift_rot_result_nxt[8]~21_combout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \R_src1[8]~23_combout ;
wire \E_src1[8]~q ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[9]~2_combout ;
wire \Add0~86 ;
wire \Add0~9_sumout ;
wire \R_src1[9]~4_combout ;
wire \E_src1[9]~q ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[10]~24_combout ;
wire \Add0~10 ;
wire \Add0~97_sumout ;
wire \R_src1[10]~26_combout ;
wire \E_src1[10]~q ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[11]~23_combout ;
wire \Add0~98 ;
wire \Add0~93_sumout ;
wire \R_src1[11]~25_combout ;
wire \E_src1[11]~q ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[12]~22_combout ;
wire \Add0~94 ;
wire \Add0~89_sumout ;
wire \R_src1[12]~24_combout ;
wire \E_src1[12]~q ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[13]~18_combout ;
wire \F_iw[17]~35_combout ;
wire \F_iw[17]~25_combout ;
wire \D_iw[17]~q ;
wire \Add0~90 ;
wire \Add0~73_sumout ;
wire \R_src1[13]~20_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[14]~17_combout ;
wire \F_iw[18]~48_combout ;
wire \F_iw[18]~26_combout ;
wire \D_iw[18]~q ;
wire \Add0~74 ;
wire \Add0~69_sumout ;
wire \R_src1[14]~19_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[15]~16_combout ;
wire \Add0~70 ;
wire \Add0~65_sumout ;
wire \F_iw[19]~63_combout ;
wire \F_iw[19]~31_combout ;
wire \D_iw[19]~q ;
wire \R_src1[15]~18_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[16]~15_combout ;
wire \Add0~66 ;
wire \Add0~61_sumout ;
wire \F_iw[20]~62_combout ;
wire \F_iw[20]~30_combout ;
wire \D_iw[20]~q ;
wire \R_src1[16]~17_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[17]~14_combout ;
wire \Add0~62 ;
wire \Add0~57_sumout ;
wire \F_iw[21]~61_combout ;
wire \F_iw[21]~21_combout ;
wire \D_iw[21]~q ;
wire \R_src1[17]~16_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[18]~13_combout ;
wire \F_iw[22]~36_combout ;
wire \F_iw[22]~0_combout ;
wire \D_iw[22]~q ;
wire \Add0~58 ;
wire \Add0~53_sumout ;
wire \R_src1[18]~15_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[19]~9_combout ;
wire \F_iw[23]~32_combout ;
wire \F_iw[23]~1_combout ;
wire \D_iw[23]~q ;
wire \Add0~54 ;
wire \Add0~37_sumout ;
wire \R_src1[19]~11_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[20]~8_combout ;
wire \F_iw[24]~37_combout ;
wire \F_iw[24]~2_combout ;
wire \D_iw[24]~q ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \R_src1[20]~10_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[21]~10_combout ;
wire \F_iw[25]~38_combout ;
wire \F_iw[25]~3_combout ;
wire \D_iw[25]~q ;
wire \Add0~34 ;
wire \Add0~41_sumout ;
wire \R_src1[21]~12_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[22]~11_combout ;
wire \F_iw[26]~39_combout ;
wire \F_iw[26]~4_combout ;
wire \D_iw[26]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \R_src1[22]~13_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[23]~12_combout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \F_iw[27]~53_combout ;
wire \F_iw[27]~27_combout ;
wire \D_iw[27]~q ;
wire \R_src1[23]~14_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[24]~3_combout ;
wire \Add0~50 ;
wire \Add0~13_sumout ;
wire \F_iw[28]~49_combout ;
wire \F_iw[28]~20_combout ;
wire \D_iw[28]~q ;
wire \R_src1[24]~5_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[25]~4_combout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \F_iw[29]~50_combout ;
wire \F_iw[29]~22_combout ;
wire \D_iw[29]~q ;
wire \R_src1[25]~6_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[26]~5_combout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \F_iw[30]~51_combout ;
wire \F_iw[30]~23_combout ;
wire \D_iw[30]~q ;
wire \R_src1[26]~7_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[27]~6_combout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \F_iw[31]~52_combout ;
wire \F_iw[31]~24_combout ;
wire \D_iw[31]~q ;
wire \R_src1[27]~8_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[28]~7_combout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \R_src1[28]~9_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[29]~27_combout ;
wire \R_src1[29]~31_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[30]~30_combout ;
wire \R_src1[30]~30_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[31]~31_combout ;
wire \R_src1[31]~29_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[0]~29_combout ;
wire \E_shift_rot_result[0]~q ;
wire \E_shift_rot_result_nxt[1]~28_combout ;
wire \R_src1[1]~32_combout ;
wire \E_src1[1]~q ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[2]~25_combout ;
wire \Add0~101_sumout ;
wire \R_src1[2]~27_combout ;
wire \E_src1[2]~q ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[3]~26_combout ;
wire \Add0~105_sumout ;
wire \R_src1[3]~28_combout ;
wire \E_src1[3]~q ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[4]~0_combout ;
wire \Add0~1_sumout ;
wire \R_src1[4]~2_combout ;
wire \E_src1[4]~q ;
wire \E_shift_rot_result[4]~q ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~0_combout ;
wire \D_ctrl_alu_force_xor~1_combout ;
wire \D_ctrl_alu_force_xor~3_combout ;
wire \D_ctrl_alu_force_xor~2_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[4]~0_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \Add2~122_cout ;
wire \Add2~114 ;
wire \Add2~110 ;
wire \Add2~102 ;
wire \Add2~106 ;
wire \Add2~1_sumout ;
wire \E_alu_result[4]~0_combout ;
wire \Equal62~3_combout ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal0~1_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;
wire \Equal62~4_combout ;
wire \Equal62~5_combout ;
wire \D_ctrl_br_cmp~0_combout ;
wire \Equal0~7_combout ;
wire \Equal0~2_combout ;
wire \Equal0~8_combout ;
wire \D_ctrl_br_cmp~1_combout ;
wire \D_ctrl_br_cmp~2_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~1_combout ;
wire \E_src2[5]~0_combout ;
wire \E_src2[5]~q ;
wire \E_logic_result[5]~1_combout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \E_alu_result[5]~2_combout ;
wire \E_src2[9]~q ;
wire \E_logic_result[9]~2_combout ;
wire \E_src2[8]~q ;
wire \E_src2[7]~q ;
wire \E_src2[6]~q ;
wire \Add2~6 ;
wire \Add2~78 ;
wire \Add2~82 ;
wire \Add2~86 ;
wire \Add2~9_sumout ;
wire \E_alu_result[9]~3_combout ;
wire \R_src2_hi[8]~0_combout ;
wire \D_ctrl_logic~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~0_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~1_combout ;
wire \E_src2[24]~q ;
wire \E_logic_result[24]~3_combout ;
wire \R_src2_hi[7]~10_combout ;
wire \E_src2[23]~q ;
wire \R_src2_hi[6]~9_combout ;
wire \E_src2[22]~q ;
wire \R_src2_hi[5]~8_combout ;
wire \E_src2[21]~q ;
wire \R_src2_hi[4]~6_combout ;
wire \E_src2[20]~q ;
wire \R_src2_hi[3]~7_combout ;
wire \E_src2[19]~q ;
wire \R_src2_hi[2]~11_combout ;
wire \E_src2[18]~q ;
wire \R_src2_hi[1]~12_combout ;
wire \E_src2[17]~q ;
wire \R_src2_hi[0]~13_combout ;
wire \E_src2[16]~q ;
wire \E_src2[15]~q ;
wire \E_src2[14]~q ;
wire \E_src2[13]~q ;
wire \E_src2[12]~q ;
wire \E_src2[11]~q ;
wire \E_src2[10]~q ;
wire \Add2~10 ;
wire \Add2~98 ;
wire \Add2~94 ;
wire \Add2~90 ;
wire \Add2~74 ;
wire \Add2~70 ;
wire \Add2~66 ;
wire \Add2~62 ;
wire \Add2~58 ;
wire \Add2~54 ;
wire \Add2~38 ;
wire \Add2~34 ;
wire \Add2~42 ;
wire \Add2~46 ;
wire \Add2~50 ;
wire \Add2~13_sumout ;
wire \E_alu_result[24]~4_combout ;
wire \R_src2_hi[9]~2_combout ;
wire \E_src2[25]~q ;
wire \E_logic_result[25]~4_combout ;
wire \Add2~14 ;
wire \Add2~17_sumout ;
wire \E_alu_result[25]~5_combout ;
wire \R_src2_hi[10]~3_combout ;
wire \E_src2[26]~q ;
wire \E_logic_result[26]~5_combout ;
wire \Add2~18 ;
wire \Add2~21_sumout ;
wire \E_alu_result[26]~6_combout ;
wire \R_src2_hi[11]~4_combout ;
wire \E_src2[27]~q ;
wire \E_logic_result[27]~6_combout ;
wire \Add2~22 ;
wire \Add2~25_sumout ;
wire \E_alu_result[27]~7_combout ;
wire \R_src2_hi[12]~5_combout ;
wire \E_src2[28]~q ;
wire \E_logic_result[28]~7_combout ;
wire \Add2~26 ;
wire \Add2~29_sumout ;
wire \E_alu_result[28]~8_combout ;
wire \E_logic_result[20]~8_combout ;
wire \Add2~33_sumout ;
wire \E_alu_result[20]~9_combout ;
wire \E_logic_result[19]~9_combout ;
wire \Add2~37_sumout ;
wire \E_alu_result[19]~10_combout ;
wire \E_logic_result[21]~10_combout ;
wire \Add2~41_sumout ;
wire \E_alu_result[21]~11_combout ;
wire \E_logic_result[22]~11_combout ;
wire \Add2~45_sumout ;
wire \E_alu_result[22]~12_combout ;
wire \E_logic_result[23]~12_combout ;
wire \Add2~49_sumout ;
wire \E_alu_result[23]~13_combout ;
wire \E_logic_result[18]~13_combout ;
wire \Add2~53_sumout ;
wire \E_alu_result[18]~14_combout ;
wire \E_logic_result[17]~14_combout ;
wire \Add2~57_sumout ;
wire \E_alu_result[17]~15_combout ;
wire \E_logic_result[16]~15_combout ;
wire \Add2~61_sumout ;
wire \E_alu_result[16]~16_combout ;
wire \E_logic_result[15]~16_combout ;
wire \Add2~65_sumout ;
wire \E_alu_result[15]~17_combout ;
wire \E_logic_result[14]~17_combout ;
wire \Add2~69_sumout ;
wire \E_alu_result[14]~18_combout ;
wire \E_logic_result[13]~18_combout ;
wire \Add2~73_sumout ;
wire \E_alu_result[13]~19_combout ;
wire \E_logic_result[6]~19_combout ;
wire \Add2~77_sumout ;
wire \E_alu_result[6]~20_combout ;
wire \E_logic_result[7]~20_combout ;
wire \Add2~81_sumout ;
wire \E_alu_result[7]~21_combout ;
wire \E_logic_result[8]~21_combout ;
wire \Add2~85_sumout ;
wire \E_alu_result[8]~22_combout ;
wire \E_logic_result[12]~22_combout ;
wire \Add2~89_sumout ;
wire \E_alu_result[12]~23_combout ;
wire \E_logic_result[11]~23_combout ;
wire \Add2~93_sumout ;
wire \E_alu_result[11]~24_combout ;
wire \E_logic_result[10]~24_combout ;
wire \Add2~97_sumout ;
wire \E_alu_result[10]~25_combout ;
wire \E_logic_result[2]~25_combout ;
wire \Add2~101_sumout ;
wire \E_alu_result[2]~26_combout ;
wire \E_logic_result[3]~26_combout ;
wire \Add2~105_sumout ;
wire \E_alu_result[3]~27_combout ;
wire \F_pc_sel_nxt.01~0_combout ;
wire \Equal0~14_combout ;
wire \Equal62~2_combout ;
wire \Equal0~3_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \R_src2_hi[15]~14_combout ;
wire \E_src2[31]~q ;
wire \R_src2_hi[14]~15_combout ;
wire \E_src2[30]~q ;
wire \R_src2_hi[13]~16_combout ;
wire \E_src2[29]~q ;
wire \Add2~30 ;
wire \Add2~134 ;
wire \Add2~130 ;
wire \Add2~126 ;
wire \Add2~117_sumout ;
wire \R_compare_op[0]~q ;
wire \E_logic_result[31]~27_combout ;
wire \E_logic_result[30]~28_combout ;
wire \E_logic_result[29]~29_combout ;
wire \E_logic_result[1]~30_combout ;
wire \E_logic_result[0]~31_combout ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \Equal127~5_combout ;
wire \Equal127~6_combout ;
wire \Equal127~7_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \Equal127~10_combout ;
wire \Equal127~11_combout ;
wire \Equal127~12_combout ;
wire \R_compare_op[1]~q ;
wire \E_cmp_result~0_combout ;
wire \W_cmp_result~q ;
wire \Equal62~11_combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~4_combout ;
wire \R_ctrl_br_uncond~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \F_pc_no_crst_nxt[17]~1_combout ;
wire \F_pc_no_crst_nxt[16]~2_combout ;
wire \F_pc_no_crst_nxt[18]~3_combout ;
wire \F_pc_no_crst_nxt[19]~4_combout ;
wire \F_pc_no_crst_nxt[20]~5_combout ;
wire \F_pc_no_crst_nxt[21]~6_combout ;
wire \F_pc_no_crst_nxt[22]~7_combout ;
wire \F_pc_no_crst_nxt[23]~8_combout ;
wire \F_pc_no_crst_nxt[24]~9_combout ;
wire \F_pc_no_crst_nxt[26]~10_combout ;
wire \F_pc_no_crst_nxt[15]~11_combout ;
wire \F_pc_no_crst_nxt[14]~12_combout ;
wire \F_pc_no_crst_nxt[9]~13_combout ;
wire \F_pc_no_crst_nxt[11]~14_combout ;
wire \F_pc_no_crst_nxt[13]~15_combout ;
wire \F_pc_no_crst_nxt[12]~16_combout ;
wire \F_pc_no_crst_nxt[10]~17_combout ;
wire \F_pc_no_crst_nxt[0]~18_combout ;
wire \F_pc_no_crst_nxt[1]~19_combout ;
wire \F_pc_no_crst_nxt[2]~20_combout ;
wire \F_pc_no_crst_nxt~21_combout ;
wire \F_pc_no_crst_nxt[4]~22_combout ;
wire \F_pc_no_crst_nxt[5]~23_combout ;
wire \F_pc_no_crst_nxt[6]~24_combout ;
wire \F_pc_no_crst_nxt[7]~25_combout ;
wire \F_pc_no_crst_nxt[8]~26_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \E_st_data[23]~0_combout ;
wire \d_read_nxt~combout ;
wire \i_read_nxt~0_combout ;
wire \F_pc_no_crst_nxt[25]~0_combout ;
wire \Add2~109_sumout ;
wire \Add2~113_sumout ;
wire \D_ctrl_mem16~1_combout ;
wire \E_mem_byte_en~0_combout ;
wire \E_mem_byte_en[1]~1_combout ;
wire \E_mem_byte_en[2]~2_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \hbreak_enabled~0_combout ;
wire \E_st_data[24]~1_combout ;
wire \E_st_data[25]~2_combout ;
wire \E_st_data[26]~3_combout ;
wire \E_st_data[27]~4_combout ;
wire \E_st_data[28]~5_combout ;
wire \E_st_data[29]~6_combout ;
wire \E_st_data[30]~7_combout ;
wire \E_st_data[31]~8_combout ;


sdram_demo_sdram_demo_nios2_cpu_register_bank_a_module sdram_demo_nios2_cpu_register_bank_a(
	.q_b_4(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_9(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.D_iw_28(\D_iw[28]~q ),
	.q_b_24(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.D_iw_29(\D_iw[29]~q ),
	.q_b_25(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.D_iw_30(\D_iw[30]~q ),
	.q_b_26(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.D_iw_31(\D_iw[31]~q ),
	.q_b_27(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_20(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_21(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_22(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.D_iw_27(\D_iw[27]~q ),
	.q_b_23(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_18(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_6(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_8(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_12(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_2(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_31(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_1(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~31_combout ),
	.W_rf_wren(\W_rf_wren~combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~0_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~1_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~2_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~3_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~4_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~5_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~6_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~7_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~8_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~9_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~10_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~11_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~12_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~13_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~14_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~15_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~16_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~17_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~18_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~19_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~20_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~21_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~22_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~23_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~24_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~25_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~26_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~27_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~28_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~29_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~30_combout ),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_nios2_oci the_sdram_demo_nios2_cpu_nios2_oci(
	.readdata_0(readdata_0),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_1(readdata_1),
	.readdata_4(readdata_4),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.readdata_11(readdata_11),
	.readdata_12(readdata_12),
	.readdata_13(readdata_13),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_16(readdata_16),
	.readdata_5(readdata_5),
	.readdata_8(readdata_8),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_28(readdata_28),
	.readdata_21(readdata_21),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.readdata_17(readdata_17),
	.readdata_18(readdata_18),
	.readdata_27(readdata_27),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.always0(always0),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled(hbreak_enabled1),
	.jtag_break(\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|jtag_break~q ),
	.WideOr1(WideOr13),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.r_early_rst(r_early_rst),
	.oci_ienable_0(\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_single_step_mode(\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.writedata_nxt({src_payload25,src_payload24,src_payload23,src_payload21,src_payload28,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload22,src_payload31,src_payload32,src_payload27,src_payload26,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,
src_payload11,src_payload19,src_payload20,src_payload18,src_payload29,src_payload30,src_payload17,src_payload10,src_payload3,src_payload4,src_payload2,src_payload}),
	.debugaccess_nxt(src_payload1),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.resetrequest(debug_reset_request),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_register_bank_b_module sdram_demo_nios2_cpu_register_bank_b(
	.q_b_0(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.D_iw_22(\D_iw[22]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_26(\D_iw[26]~q ),
	.q_b_9(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_24(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_25(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_26(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_27(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_20(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_21(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_22(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_18(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_8(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_12(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_31(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~31_combout ),
	.W_rf_wren(\W_rf_wren~combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~0_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~1_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~2_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~3_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~4_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~5_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~6_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~7_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~8_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~9_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~10_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~11_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~12_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~13_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~14_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~15_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~16_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~17_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~18_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~19_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~20_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~21_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~22_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~23_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~24_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~25_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~26_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~27_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~28_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~29_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~30_combout ),
	.clk_clk(clk_clk));

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(src_data_0),
	.asdata(\av_ld_byte1_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\E_alu_result[0]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(src_data_1),
	.asdata(\av_ld_byte1_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\E_alu_result[1]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(src_data_2),
	.asdata(\av_ld_byte1_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(src_data_3),
	.asdata(\av_ld_byte1_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(src_data_4),
	.asdata(\av_ld_byte1_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(src_data_5),
	.asdata(\av_ld_byte1_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(src_data_6),
	.asdata(\av_ld_byte1_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(src_data_7),
	.asdata(\av_ld_byte1_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(src_data_24),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(src_data_25),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(src_data_26),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(src_data_27),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(src_data_28),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cyclonev_lcell_comb \Add2~125 (
	.dataa(!\E_invert_arith_src_msb~q ),
	.datab(!\E_alu_sub~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(\Add2~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~125_sumout ),
	.cout(\Add2~126 ),
	.shareout());
defparam \Add2~125 .extended_lut = "off";
defparam \Add2~125 .lut_mask = 64'h000055AA00009966;
defparam \Add2~125 .shared_arith = "off";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(src_data_29),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(src_data_30),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(src_data_31),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

cyclonev_lcell_comb \Add2~129 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(\Add2~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~129_sumout ),
	.cout(\Add2~130 ),
	.shareout());
defparam \Add2~129 .extended_lut = "off";
defparam \Add2~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~129 .shared_arith = "off";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

cyclonev_lcell_comb \Add2~133 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~q ),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~133_sumout ),
	.cout(\Add2~134 ),
	.shareout());
defparam \Add2~133 .extended_lut = "off";
defparam \Add2~133 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~133 .shared_arith = "off";

cyclonev_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(!\Equal132~1_combout ),
	.datab(!\D_iw[8]~q ),
	.datac(!\W_bstatus_reg~q ),
	.datad(!\D_iw[6]~q ),
	.datae(!\D_iw[7]~q ),
	.dataf(!\W_ienable_reg[0]~q ),
	.datag(!\W_ipending_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_rd_data[0]~1 .extended_lut = "on";
defparam \E_control_rd_data[0]~1 .lut_mask = 64'hFBFEFBFEFBFEFBFE;
defparam \E_control_rd_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[0]~31 (
	.dataa(!\W_cmp_result~q ),
	.datab(!\av_ld_byte0_data[0]~q ),
	.datac(!\W_control_rd_data[0]~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\R_ctrl_rd_ctl_reg~q ),
	.dataf(!\R_ctrl_br_cmp~q ),
	.datag(!\W_alu_result[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[0]~31 .extended_lut = "on";
defparam \W_rf_wr_data[0]~31 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \W_rf_wr_data[0]~31 .shared_arith = "off";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cyclonev_lcell_comb W_rf_wren(
	.dataa(!r_sync_rst),
	.datab(!\R_wr_dst_reg~q ),
	.datac(!\W_valid~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam W_rf_wren.extended_lut = "off";
defparam W_rf_wren.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam W_rf_wren.shared_arith = "off";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[1]~0 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte0_data[1]~q ),
	.datae(!\W_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[1]~0 .extended_lut = "off";
defparam \W_rf_wr_data[1]~0 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[2]~1 (
	.dataa(!W_alu_result_2),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[2]~1 .extended_lut = "off";
defparam \W_rf_wr_data[2]~1 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[3]~2 (
	.dataa(!W_alu_result_3),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[3]~2 .extended_lut = "off";
defparam \W_rf_wr_data[3]~2 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[4]~3 (
	.dataa(!W_alu_result_4),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[4]~3 .extended_lut = "off";
defparam \W_rf_wr_data[4]~3 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[5]~4 (
	.dataa(!W_alu_result_5),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[5]~4 .extended_lut = "off";
defparam \W_rf_wr_data[5]~4 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[6]~5 (
	.dataa(!W_alu_result_6),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[6]~5 .extended_lut = "off";
defparam \W_rf_wr_data[6]~5 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[7]~6 (
	.dataa(!W_alu_result_7),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[7]~6 .extended_lut = "off";
defparam \W_rf_wr_data[7]~6 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[7]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\D_iw[18]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~0 .extended_lut = "off";
defparam \D_dst_regnum[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[1]~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(!\D_dst_regnum[1]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~1 .extended_lut = "off";
defparam \D_dst_regnum[1]~1 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \D_dst_regnum[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[2]~2 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\D_iw[19]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~2 .extended_lut = "off";
defparam \D_dst_regnum[2]~2 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[2]~3 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(!\D_dst_regnum[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~3 .extended_lut = "off";
defparam \D_dst_regnum[2]~3 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[3]~4 (
	.dataa(!\D_iw[25]~q ),
	.datab(!\D_iw[20]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~4 .extended_lut = "off";
defparam \D_dst_regnum[3]~4 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[3]~5 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(!\D_dst_regnum[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~5 .extended_lut = "off";
defparam \D_dst_regnum[3]~5 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[0]~6 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\D_iw[17]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~6 .extended_lut = "off";
defparam \D_dst_regnum[0]~6 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[0]~7 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(!\D_dst_regnum[0]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~7 .extended_lut = "off";
defparam \D_dst_regnum[0]~7 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[0]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[4]~8 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~8 .extended_lut = "off";
defparam \D_dst_regnum[4]~8 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[4]~9 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(!\D_dst_regnum[4]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~9 .extended_lut = "off";
defparam \D_dst_regnum[4]~9 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[4]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_wr_dst_reg~0 (
	.dataa(!\Equal0~13_combout ),
	.datab(!\R_ctrl_br_nxt~0_combout ),
	.datac(!\R_src2_use_imm~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_wr_dst_reg~0 .extended_lut = "off";
defparam \D_wr_dst_reg~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_dst_regnum[1]~1_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[3]~5_combout ),
	.datad(!\D_dst_regnum[0]~7_combout ),
	.datae(!\D_dst_regnum[4]~9_combout ),
	.dataf(!\D_wr_dst_reg~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam D_wr_dst_reg.shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld_signed~0 .extended_lut = "off";
defparam \D_ctrl_ld_signed~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \D_ctrl_ld_signed~0 .shared_arith = "off";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

cyclonev_lcell_comb \av_ld_rshift8~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\av_ld_align_cycle[1]~q ),
	.datae(!\av_ld_align_cycle[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_rshift8~0 .extended_lut = "off";
defparam \av_ld_rshift8~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \av_ld_rshift8~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte0_data[7]~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\av_ld_align_cycle[1]~q ),
	.datae(!\av_ld_align_cycle[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[7]~0 .extended_lut = "off";
defparam \av_ld_byte0_data[7]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \av_ld_byte0_data[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(!\W_status_reg_pie~q ),
	.datab(!\Equal132~0_combout ),
	.datac(!\Equal133~0_combout ),
	.datad(!\W_estatus_reg~q ),
	.datae(!\E_control_rd_data[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_rd_data[0]~0 .extended_lut = "off";
defparam \E_control_rd_data[0]~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \E_control_rd_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0]~28 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\Add2~113_sumout ),
	.datad(!\E_logic_result[0]~31_combout ),
	.datae(!\E_shift_rot_result[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0]~28 .extended_lut = "off";
defparam \E_alu_result[0]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[0]~28 .shared_arith = "off";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[9]~7 (
	.dataa(!W_alu_result_9),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[9]~7 .extended_lut = "off";
defparam \W_rf_wr_data[9]~7 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[24]~8 (
	.dataa(!W_alu_result_24),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte3_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[24]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[24]~8 .extended_lut = "off";
defparam \W_rf_wr_data[24]~8 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[24]~8 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[25]~9 (
	.dataa(!W_alu_result_25),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte3_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[25]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[25]~9 .extended_lut = "off";
defparam \W_rf_wr_data[25]~9 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[25]~9 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[26]~10 (
	.dataa(!W_alu_result_26),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte3_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[26]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[26]~10 .extended_lut = "off";
defparam \W_rf_wr_data[26]~10 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[26]~10 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[27]~11 (
	.dataa(!W_alu_result_27),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte3_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[27]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[27]~11 .extended_lut = "off";
defparam \W_rf_wr_data[27]~11 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[27]~11 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[28]~12 (
	.dataa(!W_alu_result_28),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte3_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[28]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[28]~12 .extended_lut = "off";
defparam \W_rf_wr_data[28]~12 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[28]~12 .shared_arith = "off";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[20]~13 (
	.dataa(!W_alu_result_20),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[20]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[20]~13 .extended_lut = "off";
defparam \W_rf_wr_data[20]~13 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[20]~13 .shared_arith = "off";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[19]~14 (
	.dataa(!W_alu_result_19),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[19]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[19]~14 .extended_lut = "off";
defparam \W_rf_wr_data[19]~14 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[19]~14 .shared_arith = "off";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[21]~15 (
	.dataa(!W_alu_result_21),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[21]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[21]~15 .extended_lut = "off";
defparam \W_rf_wr_data[21]~15 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[21]~15 .shared_arith = "off";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[22]~16 (
	.dataa(!W_alu_result_22),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[22]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[22]~16 .extended_lut = "off";
defparam \W_rf_wr_data[22]~16 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[22]~16 .shared_arith = "off";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[7]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[23]~17 (
	.dataa(!W_alu_result_23),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[23]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[23]~17 .extended_lut = "off";
defparam \W_rf_wr_data[23]~17 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[23]~17 .shared_arith = "off";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[18]~18 (
	.dataa(!W_alu_result_18),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[18]~18 .extended_lut = "off";
defparam \W_rf_wr_data[18]~18 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[18]~18 .shared_arith = "off";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[1]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[17]~19 (
	.dataa(!W_alu_result_17),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[17]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[17]~19 .extended_lut = "off";
defparam \W_rf_wr_data[17]~19 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[17]~19 .shared_arith = "off";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[0]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[16]~20 (
	.dataa(!W_alu_result_16),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[16]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[16]~20 .extended_lut = "off";
defparam \W_rf_wr_data[16]~20 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[16]~20 .shared_arith = "off";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[7]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[15]~21 (
	.dataa(!W_alu_result_15),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[15]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[15]~21 .extended_lut = "off";
defparam \W_rf_wr_data[15]~21 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[15]~21 .shared_arith = "off";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[14]~22 (
	.dataa(!W_alu_result_14),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[14]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[14]~22 .extended_lut = "off";
defparam \W_rf_wr_data[14]~22 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[14]~22 .shared_arith = "off";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[5]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[13]~23 (
	.dataa(!W_alu_result_13),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[13]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[13]~23 .extended_lut = "off";
defparam \W_rf_wr_data[13]~23 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[13]~23 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[8]~24 (
	.dataa(!W_alu_result_8),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[8]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[8]~24 .extended_lut = "off";
defparam \W_rf_wr_data[8]~24 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[8]~24 .shared_arith = "off";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[4]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[12]~25 (
	.dataa(!W_alu_result_12),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[12]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[12]~25 .extended_lut = "off";
defparam \W_rf_wr_data[12]~25 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[12]~25 .shared_arith = "off";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[3]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[11]~26 (
	.dataa(!W_alu_result_11),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[11]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[11]~26 .extended_lut = "off";
defparam \W_rf_wr_data[11]~26 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[11]~26 .shared_arith = "off";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[2]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[10]~27 (
	.dataa(!W_alu_result_10),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[10]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[10]~27 .extended_lut = "off";
defparam \W_rf_wr_data[10]~27 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[10]~27 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[1]~29 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[1]~q ),
	.datad(!\Add2~109_sumout ),
	.datae(!\E_logic_result[1]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[1]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[1]~29 .extended_lut = "off";
defparam \E_alu_result[1]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[1]~29 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_align_cycle[1]~q ),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[0]~0 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a40),
	.datad(!ram_block1a8),
	.datae(!\av_ld_byte1_data_nxt[0]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[0]~0 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[0]~0 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[0]~0 .shared_arith = "off";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cyclonev_lcell_comb \av_fill_bit~0 (
	.dataa(!\av_ld_byte0_data[7]~q ),
	.datab(!\D_ctrl_mem16~1_combout ),
	.datac(!\av_ld_byte1_data[7]~q ),
	.datad(!\R_ctrl_ld_signed~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_fill_bit~0 .extended_lut = "off";
defparam \av_fill_bit~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \av_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[0]~1 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[0]~q ),
	.datad(!\av_ld_byte1_data_nxt[0]~0_combout ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[0]~1 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[0]~1 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \av_ld_byte1_data_nxt[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(!\av_ld_byte0_data[7]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_en~0 .extended_lut = "off";
defparam \av_ld_byte1_data_en~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \av_ld_byte1_data_en~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[1]~2 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a41),
	.datad(!ram_block1a9),
	.datae(!\av_ld_byte1_data_nxt[1]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[1]~2 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[1]~2 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[1]~3 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[1]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[1]~3 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[1]~3 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[4]~0 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a52),
	.datad(!ram_block1a20),
	.datae(!\av_ld_byte2_data_nxt[4]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[4]~0 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[4]~0 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[4]~1 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte3_data[4]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte2_data_nxt[4]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[4]~1 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[4]~1 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte2_data_nxt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[3]~2 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a51),
	.datad(!ram_block1a19),
	.datae(!\av_ld_byte2_data_nxt[3]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[3]~2 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[3]~2 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[3]~3 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte3_data[3]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte2_data_nxt[3]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[3]~3 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[3]~3 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte2_data_nxt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[5]~4 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a53),
	.datad(!ram_block1a21),
	.datae(!\av_ld_byte2_data_nxt[5]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[5]~4 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[5]~4 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[5]~5 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!\av_ld_byte2_data_nxt[5]~4_combout ),
	.datae(!\av_ld_byte3_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[5]~5 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[5]~5 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \av_ld_byte2_data_nxt[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[6]~6 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a54),
	.datad(!ram_block1a22),
	.datae(!\av_ld_byte2_data_nxt[6]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[6]~6 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[6]~6 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[6]~7 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!\av_ld_byte2_data_nxt[6]~6_combout ),
	.datae(!\av_ld_byte3_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[6]~7 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[6]~7 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \av_ld_byte2_data_nxt[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[7]~8 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a55),
	.datad(!ram_block1a23),
	.datae(!\av_ld_byte2_data_nxt[7]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[7]~8 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[7]~8 .lut_mask = 64'hFFFFFFB8FFFFFFB8;
defparam \av_ld_byte2_data_nxt[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[7]~9 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!\av_ld_byte2_data_nxt[7]~8_combout ),
	.datae(!\av_ld_byte3_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[7]~9 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[7]~9 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \av_ld_byte2_data_nxt[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[2]~10 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a50),
	.datad(!ram_block1a18),
	.datae(!\av_ld_byte2_data_nxt[2]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[2]~10 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[2]~10 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[2]~11 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte3_data[2]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte2_data_nxt[2]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[2]~11 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[2]~11 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte2_data_nxt[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[1]~12 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a49),
	.datad(!ram_block1a17),
	.datae(!\av_ld_byte2_data_nxt[1]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[1]~12 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[1]~12 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[1]~13 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte3_data[1]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte2_data_nxt[1]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[1]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[1]~13 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[1]~13 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte2_data_nxt[1]~13 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[0]~14 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a48),
	.datad(!ram_block1a16),
	.datae(!\av_ld_byte2_data_nxt[0]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[0]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[0]~14 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[0]~14 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte2_data_nxt[0]~14 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[0]~15 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte3_data[0]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte2_data_nxt[0]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[0]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[0]~15 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[0]~15 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte2_data_nxt[0]~15 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[7]~4 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a47),
	.datad(!ram_block1a15),
	.datae(!\av_ld_byte1_data_nxt[7]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[7]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[7]~4 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[7]~4 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[7]~4 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[7]~5 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[7]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[7]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[7]~5 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[7]~5 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[7]~5 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[6]~6 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a46),
	.datad(!ram_block1a14),
	.datae(!\av_ld_byte1_data_nxt[6]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[6]~6 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[6]~6 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[6]~7 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[6]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[6]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[6]~7 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[6]~7 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[5]~8 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a45),
	.datad(!ram_block1a13),
	.datae(!\av_ld_byte1_data_nxt[5]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[5]~8 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[5]~8 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[5]~8 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[5]~9 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[5]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[5]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[5]~9 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[5]~9 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[5]~9 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[4]~10 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a44),
	.datad(!ram_block1a12),
	.datae(!\av_ld_byte1_data_nxt[4]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[4]~10 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[4]~10 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[4]~10 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[4]~11 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[4]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[4]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[4]~11 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[4]~11 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[4]~11 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[3]~12 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a43),
	.datad(!ram_block1a11),
	.datae(!\av_ld_byte1_data_nxt[3]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[3]~12 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[3]~12 .lut_mask = 64'hFFFFFFB8FFFFFFB8;
defparam \av_ld_byte1_data_nxt[3]~12 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[3]~13 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[3]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[3]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[3]~13 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[3]~13 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[3]~13 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[2]~14 (
	.dataa(!src0_valid),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a42),
	.datad(!ram_block1a10),
	.datae(!\av_ld_byte1_data_nxt[2]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[2]~14 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[2]~14 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \av_ld_byte1_data_nxt[2]~14 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[2]~15 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_ld_byte2_data[2]~q ),
	.datad(!\av_fill_bit~0_combout ),
	.datae(!\av_ld_byte1_data_nxt[2]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[2]~15 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[2]~15 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \av_ld_byte1_data_nxt[2]~15 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[31]~28 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[7]~q ),
	.datae(!\W_alu_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[31]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[31]~28 .extended_lut = "off";
defparam \W_rf_wr_data[31]~28 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[31]~28 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[30]~29 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[6]~q ),
	.datae(!\W_alu_result[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[30]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[30]~29 .extended_lut = "off";
defparam \W_rf_wr_data[30]~29 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[30]~29 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[29]~30 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[5]~q ),
	.datae(!\W_alu_result[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[29]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[29]~30 .extended_lut = "off";
defparam \W_rf_wr_data[29]~30 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[29]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31]~30 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[31]~27_combout ),
	.datad(!\Add2~125_sumout ),
	.datae(!\E_shift_rot_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31]~30 .extended_lut = "off";
defparam \E_alu_result[31]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[31]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30]~31 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[30]~28_combout ),
	.datad(!\E_shift_rot_result[30]~q ),
	.datae(!\Add2~129_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30]~31 .extended_lut = "off";
defparam \E_alu_result[30]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[30]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29]~32 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[29]~q ),
	.datad(!\E_logic_result[29]~29_combout ),
	.datae(!\Add2~133_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29]~32 .extended_lut = "off";
defparam \E_alu_result[29]~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[29]~32 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[0]~16 (
	.dataa(!src0_valid1),
	.datab(!za_data_8),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_8),
	.dataf(!av_readdata_pre_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[0]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[0]~16 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[0]~16 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[0]~16 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[4]~17 (
	.dataa(!src0_valid1),
	.datab(!za_data_12),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_12),
	.dataf(!av_readdata_pre_121),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[4]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[4]~17 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[4]~17 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[4]~17 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[3]~18 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_11),
	.datad(!za_data_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[3]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[3]~18 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[3]~18 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[3]~18 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[2]~19 (
	.dataa(!src0_valid1),
	.datab(!za_data_10),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_10),
	.dataf(!av_readdata_pre_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[2]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[2]~19 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[2]~19 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[2]~19 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[1]~20 (
	.dataa(!src0_valid1),
	.datab(!za_data_9),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_9),
	.dataf(!av_readdata_pre_91),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[1]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[1]~20 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[1]~20 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[1]~20 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[1]~16 (
	.dataa(!src0_valid1),
	.datab(!za_data_17),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_171),
	.dataf(!av_readdata_pre_17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[1]~16 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[1]~16 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[1]~16 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[0]~17 (
	.dataa(!src0_valid1),
	.datab(!za_data_16),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_161),
	.dataf(!av_readdata_pre_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[0]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[0]~17 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[0]~17 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[0]~17 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[7]~21 (
	.dataa(!src0_valid1),
	.datab(!za_data_15),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_15),
	.dataf(!av_readdata_pre_151),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[7]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[7]~21 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[7]~21 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[7]~21 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[6]~22 (
	.dataa(!src0_valid1),
	.datab(!za_data_14),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_14),
	.dataf(!av_readdata_pre_141),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[6]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[6]~22 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[6]~22 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[6]~22 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[5]~23 (
	.dataa(!src0_valid1),
	.datab(!za_data_13),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_13),
	.dataf(!av_readdata_pre_131),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[5]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[5]~23 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[5]~23 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte1_data_nxt[5]~23 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[4]~18 (
	.dataa(!src0_valid1),
	.datab(!za_data_20),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_201),
	.dataf(!av_readdata_pre_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[4]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[4]~18 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[4]~18 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[4]~18 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[3]~19 (
	.dataa(!src0_valid1),
	.datab(!za_data_19),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_191),
	.dataf(!av_readdata_pre_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[3]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[3]~19 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[3]~19 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[3]~19 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[5]~20 (
	.dataa(!src0_valid1),
	.datab(!za_data_21),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_211),
	.dataf(!av_readdata_pre_21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[5]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[5]~20 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[5]~20 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[5]~20 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[6]~21 (
	.dataa(!src0_valid1),
	.datab(!za_data_22),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_221),
	.dataf(!av_readdata_pre_22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[6]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[6]~21 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[6]~21 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[6]~21 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[7]~22 (
	.dataa(!src0_valid2),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!za_data_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[7]~22 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[7]~22 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[7]~22 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[2]~23 (
	.dataa(!src0_valid1),
	.datab(!za_data_18),
	.datac(!read_latency_shift_reg_0),
	.datad(!src0_valid2),
	.datae(!av_readdata_pre_181),
	.dataf(!av_readdata_pre_18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[2]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[2]~23 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[2]~23 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \av_ld_byte2_data_nxt[2]~23 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(!\D_iw[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 64'hFFFFFFFFBBF3FFFF;
defparam \D_ctrl_implicit_dst_eretaddr~2 .shared_arith = "off";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_24),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_25),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_26),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_27),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_28),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_20),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_19),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_21),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_22),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_23),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_18),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_17),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\E_alu_result[16]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \F_pc[17] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[17]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_17),
	.prn(vcc));
defparam \F_pc[17] .is_wysiwyg = "true";
defparam \F_pc[17] .power_up = "low";

dffeas \F_pc[16] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[16]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_16),
	.prn(vcc));
defparam \F_pc[16] .is_wysiwyg = "true";
defparam \F_pc[16] .power_up = "low";

dffeas \F_pc[18] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[18]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_18),
	.prn(vcc));
defparam \F_pc[18] .is_wysiwyg = "true";
defparam \F_pc[18] .power_up = "low";

dffeas \F_pc[19] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[19]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_19),
	.prn(vcc));
defparam \F_pc[19] .is_wysiwyg = "true";
defparam \F_pc[19] .power_up = "low";

dffeas \F_pc[20] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[20]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_20),
	.prn(vcc));
defparam \F_pc[20] .is_wysiwyg = "true";
defparam \F_pc[20] .power_up = "low";

dffeas \F_pc[21] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[21]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_21),
	.prn(vcc));
defparam \F_pc[21] .is_wysiwyg = "true";
defparam \F_pc[21] .power_up = "low";

dffeas \F_pc[22] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[22]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_22),
	.prn(vcc));
defparam \F_pc[22] .is_wysiwyg = "true";
defparam \F_pc[22] .power_up = "low";

dffeas \F_pc[23] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[23]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_23),
	.prn(vcc));
defparam \F_pc[23] .is_wysiwyg = "true";
defparam \F_pc[23] .power_up = "low";

dffeas \F_pc[24] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[24]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_24),
	.prn(vcc));
defparam \F_pc[24] .is_wysiwyg = "true";
defparam \F_pc[24] .power_up = "low";

dffeas \F_pc[26] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[26]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_26),
	.prn(vcc));
defparam \F_pc[26] .is_wysiwyg = "true";
defparam \F_pc[26] .power_up = "low";

dffeas \F_pc[15] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[15]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_15),
	.prn(vcc));
defparam \F_pc[15] .is_wysiwyg = "true";
defparam \F_pc[15] .power_up = "low";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[14]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_ctrl_exception~q ),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[25] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[25]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_25),
	.prn(vcc));
defparam \F_pc[25] .is_wysiwyg = "true";
defparam \F_pc[25] .power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

cyclonev_lcell_comb \F_iw[0]~41 (
	.dataa(!src1_valid2),
	.datab(!za_data_0),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[0]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[0]~41 .extended_lut = "off";
defparam \F_iw[0]~41 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[0]~41 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[0]~5 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!ram_block1a32),
	.datad(!address_reg_a_0),
	.datae(!ram_block1a0),
	.dataf(!\F_iw[0]~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[0]~5 .extended_lut = "off";
defparam \F_iw[0]~5 .lut_mask = 64'hAF3FFFFFFFFFFFFF;
defparam \F_iw[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \F_valid~0 (
	.dataa(!i_read1),
	.datab(!src1_valid),
	.datac(!src1_valid1),
	.datad(!src1_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_valid~0 .extended_lut = "off";
defparam \F_valid~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \F_valid~0 .shared_arith = "off";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cyclonev_lcell_comb \F_iw[1]~57 (
	.dataa(!src1_valid2),
	.datab(!za_data_1),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~57 .extended_lut = "off";
defparam \F_iw[1]~57 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[1]~57 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[1]~6 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a33),
	.datae(!ram_block1a1),
	.dataf(!\F_iw[1]~57_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~6 .extended_lut = "off";
defparam \F_iw[1]~6 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[1]~6 .shared_arith = "off";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cyclonev_lcell_comb \F_iw[4]~59 (
	.dataa(!src1_valid2),
	.datab(!za_data_4),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~59 .extended_lut = "off";
defparam \F_iw[4]~59 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[4]~59 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[4]~7 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a36),
	.datae(!ram_block1a4),
	.dataf(!\F_iw[4]~59_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~7 .extended_lut = "off";
defparam \F_iw[4]~7 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[4]~7 .shared_arith = "off";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[3]~58 (
	.dataa(!src1_valid2),
	.datab(!za_data_3),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~58 .extended_lut = "off";
defparam \F_iw[3]~58 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[3]~58 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[3]~8 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a35),
	.datae(!ram_block1a3),
	.dataf(!\F_iw[3]~58_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~8 .extended_lut = "off";
defparam \F_iw[3]~8 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[3]~8 .shared_arith = "off";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_st~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_st~0 .extended_lut = "off";
defparam \D_ctrl_st~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \D_ctrl_st~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[2]~42 (
	.dataa(!src1_valid2),
	.datab(!za_data_2),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[2]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[2]~42 .extended_lut = "off";
defparam \F_iw[2]~42 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[2]~42 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[2]~9 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a34),
	.datae(!ram_block1a2),
	.dataf(!\F_iw[2]~42_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[2]~9 .extended_lut = "off";
defparam \F_iw[2]~9 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[2]~9 .shared_arith = "off";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cyclonev_lcell_comb \d_write_nxt~0 (
	.dataa(!\E_new_inst~q ),
	.datab(!\R_ctrl_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~0 .extended_lut = "off";
defparam \d_write_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \d_write_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb E_st_stall(
	.dataa(!d_write1),
	.datab(!\d_write_nxt~0_combout ),
	.datac(!av_waitrequest),
	.datad(!sink_ready),
	.datae(!WideOr0),
	.dataf(!av_waitrequest1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_st_stall.extended_lut = "off";
defparam E_st_stall.lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam E_st_stall.shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_ld~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld~0 .extended_lut = "off";
defparam \D_ctrl_ld~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_ctrl_ld~0 .shared_arith = "off";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

cyclonev_lcell_comb \E_ld_stall~0 (
	.dataa(!\E_new_inst~q ),
	.datab(!\R_ctrl_ld~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_stall~0 .extended_lut = "off";
defparam \E_ld_stall~0 .lut_mask = 64'h7777777777777777;
defparam \E_ld_stall~0 .shared_arith = "off";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cyclonev_lcell_comb \D_ctrl_mem16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem16~0 .extended_lut = "off";
defparam \D_ctrl_mem16~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_mem16~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_align_cycle_nxt[0]~1 (
	.dataa(!d_read1),
	.datab(!WideOr11),
	.datac(!\av_ld_align_cycle[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_align_cycle_nxt[0]~1 .extended_lut = "off";
defparam \av_ld_align_cycle_nxt[0]~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \av_ld_align_cycle_nxt[0]~1 .shared_arith = "off";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cyclonev_lcell_comb \av_ld_align_cycle_nxt[1]~0 (
	.dataa(!d_read1),
	.datab(!WideOr11),
	.datac(!\av_ld_align_cycle[1]~q ),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_align_cycle_nxt[1]~0 .extended_lut = "off";
defparam \av_ld_align_cycle_nxt[1]~0 .lut_mask = 64'hBFFBBFFBBFFBBFFB;
defparam \av_ld_align_cycle_nxt[1]~0 .shared_arith = "off";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cyclonev_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(!\av_ld_align_cycle[1]~q ),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_aligning_data_nxt~0 .extended_lut = "off";
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 64'h9F6F9F6F9F6F9F6F;
defparam \av_ld_aligning_data_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem32~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem32~0 .extended_lut = "off";
defparam \D_ctrl_mem32~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_mem32~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(!d_read1),
	.datab(!WideOr11),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\av_ld_aligning_data_nxt~0_combout ),
	.datae(!\D_ctrl_mem32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_aligning_data_nxt~1 .extended_lut = "off";
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 64'hFFFFDFD5FFFFDFD5;
defparam \av_ld_aligning_data_nxt~1 .shared_arith = "off";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cyclonev_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(!d_read1),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!WideOr1),
	.datae(!\E_ld_stall~0_combout ),
	.dataf(!\av_ld_waiting_for_data~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_waiting_for_data_nxt~0 .extended_lut = "off";
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 64'hFAFFFFFFFCFFFFFF;
defparam \av_ld_waiting_for_data_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_stall~0 (
	.dataa(!\R_ctrl_ld~q ),
	.datab(!\av_ld_waiting_for_data_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~0 .extended_lut = "off";
defparam \E_stall~0 .lut_mask = 64'h7777777777777777;
defparam \E_stall~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[6]~43 (
	.dataa(!src1_valid2),
	.datab(!za_data_6),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[6]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[6]~43 .extended_lut = "off";
defparam \F_iw[6]~43 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[6]~43 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[6]~29 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a38),
	.datae(!ram_block1a6),
	.dataf(!\F_iw[6]~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[6]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[6]~29 .extended_lut = "off";
defparam \F_iw[6]~29 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[6]~29 .shared_arith = "off";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cyclonev_lcell_comb \F_iw[5]~60 (
	.dataa(!src1_valid2),
	.datab(!za_data_5),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~60 .extended_lut = "off";
defparam \F_iw[5]~60 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[5]~60 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[5]~16 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a37),
	.datae(!ram_block1a5),
	.dataf(!\F_iw[5]~60_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~16 .extended_lut = "off";
defparam \F_iw[5]~16 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[5]~16 .shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(!\D_iw[3]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[0]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(!\D_iw[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \D_ctrl_b_is_dst~0 .lut_mask = 64'hFFFF9669FFFF6996;
defparam \D_ctrl_b_is_dst~0 .shared_arith = "off";

cyclonev_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[5]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_ctrl_br_nxt~0 .extended_lut = "off";
defparam \R_ctrl_br_nxt~0 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \R_ctrl_br_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[13]~54 (
	.dataa(!src1_valid2),
	.datab(!za_data_13),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~54 .extended_lut = "off";
defparam \F_iw[13]~54 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[13]~54 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[13]~12 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a45),
	.datae(!ram_block1a13),
	.dataf(!\F_iw[13]~54_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~12 .extended_lut = "off";
defparam \F_iw[13]~12 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[13]~12 .shared_arith = "off";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cyclonev_lcell_comb \F_iw[12]~40 (
	.dataa(!src1_valid2),
	.datab(!za_data_12),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[12]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[12]~40 .extended_lut = "off";
defparam \F_iw[12]~40 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[12]~40 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[12]~11 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a44),
	.datae(!ram_block1a12),
	.dataf(!\F_iw[12]~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[12]~11 .extended_lut = "off";
defparam \F_iw[12]~11 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[12]~11 .shared_arith = "off";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cyclonev_lcell_comb \F_iw[15]~55 (
	.dataa(!src1_valid2),
	.datab(!za_data_15),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~55 .extended_lut = "off";
defparam \F_iw[15]~55 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[15]~55 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[15]~14 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a47),
	.datae(!ram_block1a15),
	.dataf(!\F_iw[15]~55_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~14 .extended_lut = "off";
defparam \F_iw[15]~14 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[15]~14 .shared_arith = "off";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

cyclonev_lcell_comb \F_iw[11]~33 (
	.dataa(!src1_valid),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_11),
	.datad(!za_data_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~33 .extended_lut = "off";
defparam \F_iw[11]~33 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[11]~33 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[11]~10 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a43),
	.datae(!ram_block1a11),
	.dataf(!\F_iw[11]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~10 .extended_lut = "off";
defparam \F_iw[11]~10 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[11]~10 .shared_arith = "off";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cyclonev_lcell_comb \F_iw[14]~34 (
	.dataa(!src1_valid2),
	.datab(!za_data_14),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[14]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[14]~34 .extended_lut = "off";
defparam \F_iw[14]~34 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[14]~34 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[14]~13 (
	.dataa(!src1_valid1),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a46),
	.datad(!ram_block1a14),
	.datae(!\intr_req~combout ),
	.dataf(!\F_iw[14]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[14]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[14]~13 .extended_lut = "off";
defparam \F_iw[14]~13 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \F_iw[14]~13 .shared_arith = "off";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cyclonev_lcell_comb \R_src2_use_imm~1 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[14]~q ),
	.dataf(!\Equal0~0_combout ),
	.datag(!\D_iw[16]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~1 .extended_lut = "on";
defparam \R_src2_use_imm~1 .lut_mask = 64'hDFFFFDFFDFFFFDFF;
defparam \R_src2_use_imm~1 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_use_imm~5 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~5 .extended_lut = "off";
defparam \R_src2_use_imm~5 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \R_src2_use_imm~5 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_use_imm~0 (
	.dataa(!\R_valid~q ),
	.datab(!\D_ctrl_b_is_dst~0_combout ),
	.datac(!\R_ctrl_br_nxt~0_combout ),
	.datad(!\R_src2_use_imm~1_combout ),
	.datae(!\R_src2_use_imm~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~0 .extended_lut = "off";
defparam \R_src2_use_imm~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \R_src2_use_imm~0 .shared_arith = "off";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cyclonev_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_src_imm5_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 64'hBBF3BBF3BBF3BBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\D_ctrl_src_imm5_shift_rot~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_src_imm5_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .shared_arith = "off";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cyclonev_lcell_comb \R_src2_lo~0 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo~0 .extended_lut = "off";
defparam \R_src2_lo~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \R_src2_lo~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \D_ctrl_hi_imm16~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \D_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cyclonev_lcell_comb \Equal62~6 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~6 .extended_lut = "off";
defparam \Equal62~6 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \Equal62~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~7 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~7 .extended_lut = "off";
defparam \Equal62~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal62~7 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~6 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~6 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~6 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \D_ctrl_implicit_dst_eretaddr~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~5 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~5 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~5 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \D_ctrl_implicit_dst_eretaddr~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~4 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~4 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~4 .lut_mask = 64'hFF69FF96FFFFFFFF;
defparam \D_ctrl_implicit_dst_eretaddr~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(!\Equal62~6_combout ),
	.datab(!\Equal62~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~12 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~12 .extended_lut = "off";
defparam \Equal0~12 .lut_mask = 64'hFFFFFBFFFFFFFFFF;
defparam \Equal0~12 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~6 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 64'h7FFFFF7FFFFFFFFF;
defparam \D_ctrl_force_src2_zero~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~5 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 64'hFFBFFFFFFFFFFFBF;
defparam \D_ctrl_force_src2_zero~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~4 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_force_src2_zero~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(!\Equal0~12_combout ),
	.datab(!\D_ctrl_force_src2_zero~6_combout ),
	.datac(!\D_ctrl_force_src2_zero~5_combout ),
	.datad(!\D_ctrl_force_src2_zero~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~0 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_force_src2_zero~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~8 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~8 .extended_lut = "off";
defparam \Equal62~8 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \Equal62~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~9 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~9 .extended_lut = "off";
defparam \Equal62~9 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \Equal62~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~10 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~10 .extended_lut = "off";
defparam \Equal62~10 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \Equal62~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~12 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~12 .extended_lut = "off";
defparam \Equal62~12 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \Equal62~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~13 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~13 .extended_lut = "off";
defparam \Equal62~13 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \Equal62~13 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(!\Equal62~8_combout ),
	.datab(!\Equal62~9_combout ),
	.datac(!\Equal62~10_combout ),
	.datad(!\Equal62~12_combout ),
	.datae(!\Equal62~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~1 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_force_src2_zero~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~9 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~9 .extended_lut = "off";
defparam \Equal0~9 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~10 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~10 .extended_lut = "off";
defparam \Equal0~10 .lut_mask = 64'hFFFFFFFFFFFFFFFB;
defparam \Equal0~10 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~2 .extended_lut = "off";
defparam \D_ctrl_retaddr~2 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \D_ctrl_retaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\Equal0~10_combout ),
	.datad(!\D_ctrl_retaddr~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~13 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~13 .extended_lut = "off";
defparam \Equal0~13 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal0~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~14 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~14 .extended_lut = "off";
defparam \Equal62~14 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal62~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~15 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~15 .extended_lut = "off";
defparam \Equal62~15 .lut_mask = 64'hFFFFFFFFFFFFFDFF;
defparam \Equal62~15 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~13_combout ),
	.datac(!\Equal62~14_combout ),
	.datad(!\Equal62~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~2 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_force_src2_zero~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datac(!\D_ctrl_force_src2_zero~0_combout ),
	.datad(!\D_ctrl_force_src2_zero~1_combout ),
	.datae(!\D_ctrl_retaddr~0_combout ),
	.dataf(!\D_ctrl_force_src2_zero~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~3 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \D_ctrl_force_src2_zero~3 .shared_arith = "off";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cyclonev_lcell_comb \R_src2_lo[0]~5 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\D_iw[6]~q ),
	.datac(!\R_src2_lo~0_combout ),
	.datad(!\R_ctrl_hi_imm16~q ),
	.datae(!\R_ctrl_force_src2_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[0]~5 .extended_lut = "off";
defparam \R_src2_lo[0]~5 .lut_mask = 64'hFF7FF777FF7FF777;
defparam \R_src2_lo[0]~5 .shared_arith = "off";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_cnt[0]~_wirecell (
	.dataa(!\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_cnt[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_cnt[0]~_wirecell .extended_lut = "off";
defparam \E_shift_rot_cnt[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \E_shift_rot_cnt[0]~_wirecell .shared_arith = "off";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_src2[0]~q ),
	.asdata(\E_shift_rot_cnt[0]~_wirecell_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add3~3 (
	.dataa(!\E_shift_rot_cnt[1]~q ),
	.datab(!\E_shift_rot_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~3 .extended_lut = "off";
defparam \Add3~3 .lut_mask = 64'h6666666666666666;
defparam \Add3~3 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[7]~45 (
	.dataa(!src1_valid2),
	.datab(!za_data_7),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[7]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[7]~45 .extended_lut = "off";
defparam \F_iw[7]~45 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[7]~45 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[7]~28 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a39),
	.datae(!ram_block1a7),
	.dataf(!\F_iw[7]~45_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[7]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[7]~28 .extended_lut = "off";
defparam \F_iw[7]~28 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[7]~28 .shared_arith = "off";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[1]~4 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[1]~4 .extended_lut = "off";
defparam \R_src2_lo[1]~4 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[1]~4 .shared_arith = "off";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\Add3~3_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add3~2 (
	.dataa(!\E_shift_rot_cnt[2]~q ),
	.datab(!\E_shift_rot_cnt[1]~q ),
	.datac(!\E_shift_rot_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~2 .extended_lut = "off";
defparam \Add3~2 .lut_mask = 64'h9696969696969696;
defparam \Add3~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[8]~44 (
	.dataa(!src1_valid2),
	.datab(!za_data_8),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[8]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[8]~44 .extended_lut = "off";
defparam \F_iw[8]~44 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[8]~44 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[8]~17 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a40),
	.datae(!ram_block1a8),
	.dataf(!\F_iw[8]~44_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[8]~17 .extended_lut = "off";
defparam \F_iw[8]~17 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[8]~17 .shared_arith = "off";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[2]~2 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\D_iw[8]~q ),
	.datad(!\R_ctrl_hi_imm16~q ),
	.datae(!\R_ctrl_force_src2_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[2]~2 .extended_lut = "off";
defparam \R_src2_lo[2]~2 .lut_mask = 64'hFF7FDF5FFF7FDF5F;
defparam \R_src2_lo[2]~2 .shared_arith = "off";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\Add3~2_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!\E_shift_rot_cnt[3]~q ),
	.datab(!\E_shift_rot_cnt[2]~q ),
	.datac(!\E_shift_rot_cnt[1]~q ),
	.datad(!\E_shift_rot_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h6996699669966996;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[9]~46 (
	.dataa(!src1_valid2),
	.datab(!za_data_9),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[9]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[9]~46 .extended_lut = "off";
defparam \F_iw[9]~46 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[9]~46 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[9]~19 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a41),
	.datae(!ram_block1a9),
	.dataf(!\F_iw[9]~46_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[9]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[9]~19 .extended_lut = "off";
defparam \F_iw[9]~19 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[9]~19 .shared_arith = "off";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[3]~3 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[3]~3 .extended_lut = "off";
defparam \R_src2_lo[3]~3 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[3]~3 .shared_arith = "off";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\Add3~1_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cyclonev_lcell_comb \E_stall~1 (
	.dataa(!\E_shift_rot_cnt[3]~q ),
	.datab(!\E_shift_rot_cnt[2]~q ),
	.datac(!\E_shift_rot_cnt[1]~q ),
	.datad(!\E_shift_rot_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~1 .extended_lut = "off";
defparam \E_stall~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \E_stall~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!\E_shift_rot_cnt[4]~q ),
	.datab(!\E_stall~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h6666666666666666;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[10]~47 (
	.dataa(!src1_valid2),
	.datab(!za_data_10),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[10]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[10]~47 .extended_lut = "off";
defparam \F_iw[10]~47 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[10]~47 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[10]~18 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a42),
	.datae(!ram_block1a10),
	.dataf(!\F_iw[10]~47_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[10]~18 .extended_lut = "off";
defparam \F_iw[10]~18 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[10]~18 .shared_arith = "off";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[4]~1 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[4]~1 .extended_lut = "off";
defparam \R_src2_lo[4]~1 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[4]~1 .shared_arith = "off";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\Add3~0_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cyclonev_lcell_comb \E_stall~2 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\E_new_inst~q ),
	.datac(!\E_shift_rot_cnt[4]~q ),
	.datad(!\E_stall~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~2 .extended_lut = "off";
defparam \E_stall~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_stall~2 .shared_arith = "off";

cyclonev_lcell_comb \E_stall~3 (
	.dataa(!\R_ctrl_ld~q ),
	.datab(!\D_ctrl_mem32~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~3 .extended_lut = "off";
defparam \E_stall~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \E_stall~3 .shared_arith = "off";

cyclonev_lcell_comb \E_stall~4 (
	.dataa(!\E_ld_stall~0_combout ),
	.datab(!\E_valid_from_R~q ),
	.datac(!\av_ld_aligning_data_nxt~1_combout ),
	.datad(!\E_stall~0_combout ),
	.datae(!\E_stall~2_combout ),
	.dataf(!\E_stall~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~4 .extended_lut = "off";
defparam \E_stall~4 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \E_stall~4 .shared_arith = "off";

cyclonev_lcell_comb \E_valid_from_R~0 (
	.dataa(!\E_st_stall~combout ),
	.datab(!\R_valid~q ),
	.datac(!\E_stall~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid_from_R~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid_from_R~0 .extended_lut = "off";
defparam \E_valid_from_R~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \E_valid_from_R~0 .shared_arith = "off";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cyclonev_lcell_comb \W_valid~0 (
	.dataa(!\E_st_stall~combout ),
	.datab(!\E_valid_from_R~q ),
	.datac(!\E_stall~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_valid~0 .extended_lut = "off";
defparam \W_valid~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \W_valid~0 .shared_arith = "off";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cyclonev_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\hbreak_pending~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_pending_nxt~0 .extended_lut = "off";
defparam \hbreak_pending_nxt~0 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \hbreak_pending_nxt~0 .shared_arith = "off";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\wait_for_one_post_bret_inst~q ),
	.datac(!\F_valid~0_combout ),
	.datad(!\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!\W_valid~q ),
	.datab(!hbreak_enabled1),
	.datac(!\hbreak_pending~q ),
	.datad(!\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_oci_debug|jtag_break~q ),
	.datae(!\wait_for_one_post_bret_inst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \hbreak_req~0 .shared_arith = "off";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~3 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~3 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_implicit_dst_eretaddr~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~11 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~11 .extended_lut = "off";
defparam \Equal0~11 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \Equal0~11 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\Equal0~10_combout ),
	.datab(!\Equal0~11_combout ),
	.datac(!\Equal0~12_combout ),
	.datad(!\D_ctrl_force_src2_zero~6_combout ),
	.datae(!\D_ctrl_force_src2_zero~5_combout ),
	.dataf(!\D_ctrl_force_src2_zero~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(!\D_iw[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~1 .extended_lut = "off";
defparam \D_ctrl_exception~1 .lut_mask = 64'hF7FFFFFFB3FFFFFF;
defparam \D_ctrl_exception~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.datad(!\D_ctrl_exception~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~0 .extended_lut = "off";
defparam \D_ctrl_exception~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_exception~0 .shared_arith = "off";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cyclonev_lcell_comb \D_ctrl_break~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~0 .extended_lut = "off";
defparam \D_ctrl_break~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_break~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_break~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_ctrl_break~0_combout ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~1 .extended_lut = "off";
defparam \D_ctrl_break~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \D_ctrl_break~1 .shared_arith = "off";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cyclonev_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~3 .extended_lut = "off";
defparam \D_ctrl_retaddr~3 .lut_mask = 64'hF7FFD5FFFFFFFFFF;
defparam \D_ctrl_retaddr~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datac(!\Equal0~11_combout ),
	.datad(!\D_ctrl_force_src2_zero~0_combout ),
	.datae(!\D_ctrl_retaddr~3_combout ),
	.dataf(!\D_ctrl_retaddr~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \R_src1~0 (
	.dataa(!\E_valid_from_R~q ),
	.datab(!\R_ctrl_br~q ),
	.datac(!\R_valid~q ),
	.datad(!\R_ctrl_retaddr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1~0 .extended_lut = "off";
defparam \R_src1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \R_src1~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_jmp_direct~0 .extended_lut = "off";
defparam \D_ctrl_jmp_direct~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_jmp_direct~0 .shared_arith = "off";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

cyclonev_lcell_comb \R_src1~1 (
	.dataa(!\E_valid_from_R~q ),
	.datab(!\R_ctrl_jmp_direct~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1~1 .extended_lut = "off";
defparam \R_src1~1 .lut_mask = 64'h7777777777777777;
defparam \R_src1~1 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[0]~33 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[0]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[0]~33 .extended_lut = "off";
defparam \R_src1[0]~33 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \R_src1[0]~33 .shared_arith = "off";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\R_src1[0]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cyclonev_lcell_comb \Equal132~1 (
	.dataa(!\D_iw[9]~q ),
	.datab(!\D_iw[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal132~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal132~1 .extended_lut = "off";
defparam \Equal132~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal132~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal133~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\Equal132~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal133~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal133~0 .extended_lut = "off";
defparam \Equal133~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \Equal133~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~16 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~16 .extended_lut = "off";
defparam \Equal62~16 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \Equal62~16 .shared_arith = "off";

cyclonev_lcell_comb D_op_wrctl(
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_op_wrctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_op_wrctl.extended_lut = "off";
defparam D_op_wrctl.lut_mask = 64'h7777777777777777;
defparam D_op_wrctl.shared_arith = "off";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\Equal133~0_combout ),
	.datac(!\W_estatus_reg~q ),
	.datad(!\R_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_estatus_reg_inst_nxt~0 .extended_lut = "off";
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \W_estatus_reg_inst_nxt~0 .shared_arith = "off";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~0_combout ),
	.asdata(\W_status_reg_pie~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_ctrl_exception~q ),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cyclonev_lcell_comb \Equal134~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\Equal132~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal134~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal134~0 .extended_lut = "off";
defparam \Equal134~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \Equal134~0 .shared_arith = "off";

cyclonev_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(!\W_status_reg_pie~q ),
	.datad(!\W_bstatus_reg~q ),
	.datae(!\Equal134~0_combout ),
	.dataf(!\R_ctrl_wrctl_inst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_bstatus_reg_inst_nxt~0 .extended_lut = "off";
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 64'hDFFF7FFF7FFFDFFF;
defparam \W_bstatus_reg_inst_nxt~0 .shared_arith = "off";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cyclonev_lcell_comb \Equal132~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\D_iw[9]~q ),
	.datae(!\D_iw[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal132~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal132~0 .extended_lut = "off";
defparam \Equal132~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal132~0 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\W_status_reg_pie~q ),
	.datac(!\Equal132~0_combout ),
	.datad(!\R_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \W_status_reg_pie_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\W_estatus_reg~q ),
	.datac(!\W_bstatus_reg~q ),
	.datad(!\Equal62~14_combout ),
	.datae(!\Equal62~15_combout ),
	.dataf(!\W_status_reg_pie_inst_nxt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~1 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 64'hBF7F7FBFFFFFFFFF;
defparam \W_status_reg_pie_inst_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(!\R_ctrl_exception~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(!\W_status_reg_pie_inst_nxt~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~2 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \W_status_reg_pie_inst_nxt~2 .shared_arith = "off";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cyclonev_lcell_comb \Equal135~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\Equal132~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal135~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal135~0 .extended_lut = "off";
defparam \Equal135~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Equal135~0 .shared_arith = "off";

cyclonev_lcell_comb \W_ienable_reg[0]~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\E_valid_from_R~q ),
	.datac(!\W_ienable_reg[0]~q ),
	.datad(!\Equal135~0_combout ),
	.datae(!\R_ctrl_wrctl_inst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_ienable_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_ienable_reg[0]~0 .extended_lut = "off";
defparam \W_ienable_reg[0]~0 .lut_mask = 64'hDF7F7FDFDF7F7FDF;
defparam \W_ienable_reg[0]~0 .shared_arith = "off";

dffeas \W_ienable_reg[0] (
	.clk(clk_clk),
	.d(\W_ienable_reg[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ienable_reg[0]~q ),
	.prn(vcc));
defparam \W_ienable_reg[0] .is_wysiwyg = "true";
defparam \W_ienable_reg[0] .power_up = "low";

cyclonev_lcell_comb \W_ipending_reg_nxt[0]~0 (
	.dataa(!\W_ienable_reg[0]~q ),
	.datab(!\the_sdram_demo_nios2_cpu_nios2_oci|the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.datac(!av_readdata_9),
	.datad(!av_readdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_ipending_reg_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_ipending_reg_nxt[0]~0 .extended_lut = "off";
defparam \W_ipending_reg_nxt[0]~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \W_ipending_reg_nxt[0]~0 .shared_arith = "off";

dffeas \W_ipending_reg[0] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[0]~q ),
	.prn(vcc));
defparam \W_ipending_reg[0] .is_wysiwyg = "true";
defparam \W_ipending_reg[0] .power_up = "low";

cyclonev_lcell_comb intr_req(
	.dataa(!\W_status_reg_pie~q ),
	.datab(!\W_ipending_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\intr_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam intr_req.extended_lut = "off";
defparam intr_req.lut_mask = 64'h7777777777777777;
defparam intr_req.shared_arith = "off";

cyclonev_lcell_comb \D_iw[1]~0 (
	.dataa(!\intr_req~combout ),
	.datab(!\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_iw[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_iw[1]~0 .extended_lut = "off";
defparam \D_iw[1]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \D_iw[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[16]~56 (
	.dataa(!src1_valid2),
	.datab(!za_data_16),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~56 .extended_lut = "off";
defparam \F_iw[16]~56 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[16]~56 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[16]~15 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a48),
	.datae(!ram_block1a16),
	.dataf(!\F_iw[16]~56_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~15 .extended_lut = "off";
defparam \F_iw[16]~15 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[16]~15 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot~0 .lut_mask = 64'hBFB3FFFFFFFFFFFF;
defparam \D_ctrl_shift_rot~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(gnd),
	.datab(!\D_ctrl_shift_rot~0_combout ),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot~1 .lut_mask = 64'h33FF33FF33FF33FF;
defparam \D_ctrl_shift_rot~1 .shared_arith = "off";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(!\D_ctrl_logic~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_shift_rot_right~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\D_ctrl_shift_rot_right~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_ctrl_shift_rot_right~1 .shared_arith = "off";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \Equal62~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~0 .extended_lut = "off";
defparam \Equal62~0 .lut_mask = 64'hFFFFFFFFFBFFFFFF;
defparam \Equal62~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\D_iw[13]~q ),
	.dataf(!\D_iw[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~2 .extended_lut = "off";
defparam \D_ctrl_shift_rot~2 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \D_ctrl_shift_rot~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(!\Equal62~0_combout ),
	.datab(!\D_ctrl_shift_rot~2_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_logical~0 .extended_lut = "off";
defparam \D_ctrl_shift_logical~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_shift_logical~0 .shared_arith = "off";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cyclonev_lcell_comb \Equal62~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~1 .extended_lut = "off";
defparam \Equal62~1 .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \Equal62~1 .shared_arith = "off";

cyclonev_lcell_comb R_ctrl_rot_right_nxt(
	.dataa(!\Equal62~1_combout ),
	.datab(!\Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_rot_right_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam R_ctrl_rot_right_nxt.extended_lut = "off";
defparam R_ctrl_rot_right_nxt.lut_mask = 64'h7777777777777777;
defparam R_ctrl_rot_right_nxt.shared_arith = "off";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[5]~1 (
	.dataa(!\E_shift_rot_result[4]~q ),
	.datab(!\E_shift_rot_result[6]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[5]~1 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[5]~1 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h00000000000000FF;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h00000000000000FF;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[5]~3 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[9]~q ),
	.datad(!\Add0~5_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[5]~3 .extended_lut = "off";
defparam \R_src1[5]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[5]~3 .shared_arith = "off";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\R_src1[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~1_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[6]~19 (
	.dataa(!\E_shift_rot_result[5]~q ),
	.datab(!\E_shift_rot_result[7]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[6]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[6]~19 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[6]~19 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[6]~19 .shared_arith = "off";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h00000000000000FF;
defparam \Add0~77 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[6]~21 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[10]~q ),
	.datad(!\Add0~77_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[6]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[6]~21 .extended_lut = "off";
defparam \R_src1[6]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[6]~21 .shared_arith = "off";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\R_src1[6]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~19_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[7]~20 (
	.dataa(!\E_shift_rot_result[6]~q ),
	.datab(!\E_shift_rot_result[8]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[7]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[7]~20 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[7]~20 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h00000000000000FF;
defparam \Add0~81 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[7]~22 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~81_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[7]~22 .extended_lut = "off";
defparam \R_src1[7]~22 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[7]~22 .shared_arith = "off";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\R_src1[7]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~20_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[8]~21 (
	.dataa(!\E_shift_rot_result[7]~q ),
	.datab(!\E_shift_rot_result[9]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[8]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[8]~21 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[8]~21 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[8]~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h00000000000000FF;
defparam \Add0~85 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[8]~23 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~85_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[8]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[8]~23 .extended_lut = "off";
defparam \R_src1[8]~23 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[8]~23 .shared_arith = "off";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\R_src1[8]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~21_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[9]~2 (
	.dataa(!\E_shift_rot_result[8]~q ),
	.datab(!\E_shift_rot_result[10]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[9]~2 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[9]~2 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[9]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[9]~4 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~9_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[9]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[9]~4 .extended_lut = "off";
defparam \R_src1[9]~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[9]~4 .shared_arith = "off";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\R_src1[9]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~2_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[10]~24 (
	.dataa(!\E_shift_rot_result[11]~q ),
	.datab(!\E_shift_rot_result[9]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[10]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[10]~24 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[10]~24 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[10]~24 .shared_arith = "off";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h00000000000000FF;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[10]~26 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~97_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[10]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[10]~26 .extended_lut = "off";
defparam \R_src1[10]~26 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[10]~26 .shared_arith = "off";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\R_src1[10]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~24_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[11]~23 (
	.dataa(!\E_shift_rot_result[12]~q ),
	.datab(!\E_shift_rot_result[10]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[11]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[11]~23 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[11]~23 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[11]~23 .shared_arith = "off";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h00000000000000FF;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[11]~25 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~93_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[11]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[11]~25 .extended_lut = "off";
defparam \R_src1[11]~25 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[11]~25 .shared_arith = "off";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\R_src1[11]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~23_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[12]~22 (
	.dataa(!\E_shift_rot_result[11]~q ),
	.datab(!\E_shift_rot_result[13]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[12]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[12]~22 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[12]~22 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[12]~22 .shared_arith = "off";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h00000000000000FF;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[12]~24 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~89_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[12]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[12]~24 .extended_lut = "off";
defparam \R_src1[12]~24 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[12]~24 .shared_arith = "off";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\R_src1[12]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~22_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[13]~18 (
	.dataa(!\E_shift_rot_result[12]~q ),
	.datab(!\E_shift_rot_result[14]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[13]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[13]~18 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[13]~18 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[13]~18 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[17]~35 (
	.dataa(!src1_valid2),
	.datab(!za_data_17),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[17]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[17]~35 .extended_lut = "off";
defparam \F_iw[17]~35 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[17]~35 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[17]~25 (
	.dataa(!src1_valid1),
	.datab(!address_reg_a_0),
	.datac(!ram_block1a49),
	.datad(!ram_block1a17),
	.datae(!\intr_req~combout ),
	.dataf(!\F_iw[17]~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[17]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[17]~25 .extended_lut = "off";
defparam \F_iw[17]~25 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \F_iw[17]~25 .shared_arith = "off";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h00000000000000FF;
defparam \Add0~73 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[13]~20 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[17]~q ),
	.datad(!\Add0~73_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[13]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[13]~20 .extended_lut = "off";
defparam \R_src1[13]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[13]~20 .shared_arith = "off";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\R_src1[13]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~18_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[14]~17 (
	.dataa(!\E_shift_rot_result[15]~q ),
	.datab(!\E_shift_rot_result[13]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[14]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[14]~17 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[14]~17 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[14]~17 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[18]~48 (
	.dataa(!src1_valid2),
	.datab(!\intr_req~combout ),
	.datac(!\hbreak_req~0_combout ),
	.datad(!za_data_18),
	.datae(!src1_valid),
	.dataf(!av_readdata_pre_181),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~48 .extended_lut = "off";
defparam \F_iw[18]~48 .lut_mask = 64'hFFFFFFFFFFFFFFFB;
defparam \F_iw[18]~48 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[18]~26 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a50),
	.datae(!ram_block1a18),
	.dataf(!\F_iw[18]~48_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~26 .extended_lut = "off";
defparam \F_iw[18]~26 .lut_mask = 64'hBFFFFFFFB3FFFFFF;
defparam \F_iw[18]~26 .shared_arith = "off";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[14]~19 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[18]~q ),
	.datad(!\Add0~69_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[14]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[14]~19 .extended_lut = "off";
defparam \R_src1[14]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[14]~19 .shared_arith = "off";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\R_src1[14]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~17_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[15]~16 (
	.dataa(!\E_shift_rot_result[16]~q ),
	.datab(!\E_shift_rot_result[14]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[15]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[15]~16 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[15]~16 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[15]~16 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[19]~63 (
	.dataa(!src1_valid2),
	.datab(!za_data_19),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~63 .extended_lut = "off";
defparam \F_iw[19]~63 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[19]~63 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[19]~31 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a51),
	.datae(!ram_block1a19),
	.dataf(!\F_iw[19]~63_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~31 .extended_lut = "off";
defparam \F_iw[19]~31 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[19]~31 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cyclonev_lcell_comb \R_src1[15]~18 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~65_sumout ),
	.datad(!\D_iw[19]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[15]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[15]~18 .extended_lut = "off";
defparam \R_src1[15]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[15]~18 .shared_arith = "off";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\R_src1[15]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~16_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[16]~15 (
	.dataa(!\E_shift_rot_result[17]~q ),
	.datab(!\E_shift_rot_result[15]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[16]~15 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[16]~15 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[16]~15 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[20]~62 (
	.dataa(!src1_valid2),
	.datab(!za_data_20),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~62 .extended_lut = "off";
defparam \F_iw[20]~62 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[20]~62 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[20]~30 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a52),
	.datae(!ram_block1a20),
	.dataf(!\F_iw[20]~62_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~30 .extended_lut = "off";
defparam \F_iw[20]~30 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[20]~30 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \R_src1[16]~17 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~61_sumout ),
	.datad(!\D_iw[20]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[16]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[16]~17 .extended_lut = "off";
defparam \R_src1[16]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[16]~17 .shared_arith = "off";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\R_src1[16]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~15_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[17]~14 (
	.dataa(!\E_shift_rot_result[16]~q ),
	.datab(!\E_shift_rot_result[18]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[17]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[17]~14 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[17]~14 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[17]~14 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[21]~61 (
	.dataa(!src1_valid2),
	.datab(!za_data_21),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~61 .extended_lut = "off";
defparam \F_iw[21]~61 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[21]~61 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[21]~21 (
	.dataa(!\D_iw[1]~0_combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a53),
	.datae(!ram_block1a21),
	.dataf(!\F_iw[21]~61_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~21 .extended_lut = "off";
defparam \F_iw[21]~21 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[21]~21 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclonev_lcell_comb \R_src1[17]~16 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~57_sumout ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[17]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[17]~16 .extended_lut = "off";
defparam \R_src1[17]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[17]~16 .shared_arith = "off";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\R_src1[17]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~14_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[18]~13 (
	.dataa(!\E_shift_rot_result[17]~q ),
	.datab(!\E_shift_rot_result[19]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[18]~13 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[18]~13 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[18]~13 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[22]~36 (
	.dataa(!src1_valid2),
	.datab(!za_data_22),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[22]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[22]~36 .extended_lut = "off";
defparam \F_iw[22]~36 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[22]~36 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[22]~0 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a54),
	.datae(!ram_block1a22),
	.dataf(!\F_iw[22]~36_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[22]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[22]~0 .extended_lut = "off";
defparam \F_iw[22]~0 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[22]~0 .shared_arith = "off";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[18]~15 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~53_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[18]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[18]~15 .extended_lut = "off";
defparam \R_src1[18]~15 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[18]~15 .shared_arith = "off";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\R_src1[18]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~13_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[19]~9 (
	.dataa(!\E_shift_rot_result[20]~q ),
	.datab(!\E_shift_rot_result[18]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[19]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[19]~9 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[19]~9 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[19]~9 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[23]~32 (
	.dataa(!src1_valid2),
	.datab(!za_data_23),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[23]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[23]~32 .extended_lut = "off";
defparam \F_iw[23]~32 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[23]~32 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[23]~1 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a55),
	.datae(!ram_block1a23),
	.dataf(!\F_iw[23]~32_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[23]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[23]~1 .extended_lut = "off";
defparam \F_iw[23]~1 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[23]~1 .shared_arith = "off";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[19]~11 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~37_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[19]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[19]~11 .extended_lut = "off";
defparam \R_src1[19]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[19]~11 .shared_arith = "off";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\R_src1[19]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~9_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[20]~8 (
	.dataa(!\E_shift_rot_result[19]~q ),
	.datab(!\E_shift_rot_result[21]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[20]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[20]~8 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[20]~8 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[20]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[24]~37 (
	.dataa(!src1_valid2),
	.datab(!za_data_24),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[24]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[24]~37 .extended_lut = "off";
defparam \F_iw[24]~37 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[24]~37 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[24]~2 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a56),
	.datae(!ram_block1a24),
	.dataf(!\F_iw[24]~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[24]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[24]~2 .extended_lut = "off";
defparam \F_iw[24]~2 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[24]~2 .shared_arith = "off";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[20]~10 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~33_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[20]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[20]~10 .extended_lut = "off";
defparam \R_src1[20]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[20]~10 .shared_arith = "off";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\R_src1[20]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~8_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[21]~10 (
	.dataa(!\E_shift_rot_result[20]~q ),
	.datab(!\E_shift_rot_result[22]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[21]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[21]~10 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[21]~10 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[21]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[25]~38 (
	.dataa(!src1_valid2),
	.datab(!za_data_25),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[25]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[25]~38 .extended_lut = "off";
defparam \F_iw[25]~38 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[25]~38 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[25]~3 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a57),
	.datae(!ram_block1a25),
	.dataf(!\F_iw[25]~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[25]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[25]~3 .extended_lut = "off";
defparam \F_iw[25]~3 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[25]~3 .shared_arith = "off";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[21]~12 (
	.dataa(!\D_iw[25]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~41_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[21]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[21]~12 .extended_lut = "off";
defparam \R_src1[21]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[21]~12 .shared_arith = "off";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\R_src1[21]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~10_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[22]~11 (
	.dataa(!\E_shift_rot_result[21]~q ),
	.datab(!\E_shift_rot_result[23]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[22]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[22]~11 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[22]~11 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[22]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[26]~39 (
	.dataa(!src1_valid2),
	.datab(!za_data_26),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[26]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[26]~39 .extended_lut = "off";
defparam \F_iw[26]~39 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[26]~39 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[26]~4 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a58),
	.datae(!ram_block1a26),
	.dataf(!\F_iw[26]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[26]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[26]~4 .extended_lut = "off";
defparam \F_iw[26]~4 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[26]~4 .shared_arith = "off";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[22]~13 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~45_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[22]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[22]~13 .extended_lut = "off";
defparam \R_src1[22]~13 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[22]~13 .shared_arith = "off";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\R_src1[22]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~11_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[23]~12 (
	.dataa(!\E_shift_rot_result[24]~q ),
	.datab(!\E_shift_rot_result[22]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[23]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[23]~12 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[23]~12 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[23]~12 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[27]~53 (
	.dataa(!src1_valid2),
	.datab(!za_data_27),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[27]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[27]~53 .extended_lut = "off";
defparam \F_iw[27]~53 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[27]~53 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[27]~27 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a59),
	.datae(!ram_block1a27),
	.dataf(!\F_iw[27]~53_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[27]~27 .extended_lut = "off";
defparam \F_iw[27]~27 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[27]~27 .shared_arith = "off";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cyclonev_lcell_comb \R_src1[23]~14 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~49_sumout ),
	.datad(!\D_iw[27]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[23]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[23]~14 .extended_lut = "off";
defparam \R_src1[23]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[23]~14 .shared_arith = "off";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\R_src1[23]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~12_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[24]~3 (
	.dataa(!\E_shift_rot_result[25]~q ),
	.datab(!\E_shift_rot_result[23]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[24]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[24]~3 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[24]~3 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[24]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[28]~49 (
	.dataa(!src1_valid2),
	.datab(!za_data_28),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[28]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[28]~49 .extended_lut = "off";
defparam \F_iw[28]~49 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[28]~49 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[28]~20 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a60),
	.datae(!ram_block1a28),
	.dataf(!\F_iw[28]~49_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[28]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[28]~20 .extended_lut = "off";
defparam \F_iw[28]~20 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[28]~20 .shared_arith = "off";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cyclonev_lcell_comb \R_src1[24]~5 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~13_sumout ),
	.datad(!\D_iw[28]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[24]~5 .extended_lut = "off";
defparam \R_src1[24]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[24]~5 .shared_arith = "off";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\R_src1[24]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~3_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[25]~4 (
	.dataa(!\E_shift_rot_result[24]~q ),
	.datab(!\E_shift_rot_result[26]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[25]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[25]~4 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[25]~4 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[25]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[29]~50 (
	.dataa(!src1_valid2),
	.datab(!za_data_29),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[29]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[29]~50 .extended_lut = "off";
defparam \F_iw[29]~50 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[29]~50 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[29]~22 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a61),
	.datae(!ram_block1a29),
	.dataf(!\F_iw[29]~50_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[29]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[29]~22 .extended_lut = "off";
defparam \F_iw[29]~22 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[29]~22 .shared_arith = "off";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cyclonev_lcell_comb \R_src1[25]~6 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~17_sumout ),
	.datad(!\D_iw[29]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[25]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[25]~6 .extended_lut = "off";
defparam \R_src1[25]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[25]~6 .shared_arith = "off";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\R_src1[25]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~4_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[26]~5 (
	.dataa(!\E_shift_rot_result[25]~q ),
	.datab(!\E_shift_rot_result[27]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[26]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[26]~5 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[26]~5 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[26]~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[30]~51 (
	.dataa(!src1_valid2),
	.datab(!za_data_30),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[30]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[30]~51 .extended_lut = "off";
defparam \F_iw[30]~51 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[30]~51 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[30]~23 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a62),
	.datae(!ram_block1a30),
	.dataf(!\F_iw[30]~51_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[30]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[30]~23 .extended_lut = "off";
defparam \F_iw[30]~23 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[30]~23 .shared_arith = "off";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cyclonev_lcell_comb \R_src1[26]~7 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\D_iw[30]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[26]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[26]~7 .extended_lut = "off";
defparam \R_src1[26]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[26]~7 .shared_arith = "off";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\R_src1[26]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~5_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[27]~6 (
	.dataa(!\E_shift_rot_result[26]~q ),
	.datab(!\E_shift_rot_result[28]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[27]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[27]~6 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[27]~6 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[27]~6 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[31]~52 (
	.dataa(!src1_valid2),
	.datab(!za_data_31),
	.datac(!src1_valid),
	.datad(!av_readdata_pre_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[31]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[31]~52 .extended_lut = "off";
defparam \F_iw[31]~52 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \F_iw[31]~52 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[31]~24 (
	.dataa(!\intr_req~combout ),
	.datab(!src1_valid1),
	.datac(!address_reg_a_0),
	.datad(!ram_block1a63),
	.datae(!ram_block1a31),
	.dataf(!\F_iw[31]~52_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[31]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[31]~24 .extended_lut = "off";
defparam \F_iw[31]~24 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \F_iw[31]~24 .shared_arith = "off";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cyclonev_lcell_comb \R_src1[27]~8 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~25_sumout ),
	.datad(!\D_iw[31]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[27]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[27]~8 .extended_lut = "off";
defparam \R_src1[27]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[27]~8 .shared_arith = "off";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\R_src1[27]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~6_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[28]~7 (
	.dataa(!\E_shift_rot_result[27]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[28]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[28]~7 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[28]~7 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[28]~7 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[28]~9 (
	.dataa(!F_pc_26),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~29_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[28]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[28]~9 .extended_lut = "off";
defparam \R_src1[28]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[28]~9 .shared_arith = "off";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\R_src1[28]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~7_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[29]~27 (
	.dataa(!\E_shift_rot_result[28]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[29]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[29]~27 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[29]~27 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[29]~27 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[29]~31 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[29]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[29]~31 .extended_lut = "off";
defparam \R_src1[29]~31 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \R_src1[29]~31 .shared_arith = "off";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\R_src1[29]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~27_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[30]~30 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[29]~q ),
	.datac(!\E_shift_rot_result[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[30]~30 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[30]~30 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[30]~30 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[30]~30 .extended_lut = "off";
defparam \R_src1[30]~30 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \R_src1[30]~30 .shared_arith = "off";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\R_src1[30]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~30_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[31]~31 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[30]~q ),
	.datac(!\E_shift_rot_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[31]~31 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[31]~31 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[31]~31 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[31]~29 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[31]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[31]~29 .extended_lut = "off";
defparam \R_src1[31]~29 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \R_src1[31]~29 .shared_arith = "off";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\R_src1[31]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~31_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(!\E_shift_rot_result[0]~q ),
	.datab(!\R_ctrl_shift_logical~q ),
	.datac(!\R_ctrl_rot_right~q ),
	.datad(!\E_shift_rot_result[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_fill_bit~0 .extended_lut = "off";
defparam \E_shift_rot_fill_bit~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \E_shift_rot_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \E_shift_rot_result_nxt[0]~29 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[1]~q ),
	.datac(!\E_shift_rot_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[0]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[0]~29 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[0]~29 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[0]~29 .shared_arith = "off";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~29_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[1]~28 (
	.dataa(!\E_shift_rot_result[2]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[1]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[1]~28 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[1]~28 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[1]~28 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[1]~32 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[1]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[1]~32 .extended_lut = "off";
defparam \R_src1[1]~32 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \R_src1[1]~32 .shared_arith = "off";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\R_src1[1]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~28_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[2]~25 (
	.dataa(!\E_shift_rot_result[3]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[2]~25 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[2]~25 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[2]~25 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[2]~27 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\Add0~101_sumout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\D_iw[6]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[2]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[2]~27 .extended_lut = "off";
defparam \R_src1[2]~27 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \R_src1[2]~27 .shared_arith = "off";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\R_src1[2]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~25_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[3]~26 (
	.dataa(!\E_shift_rot_result[2]~q ),
	.datab(!\E_shift_rot_result[4]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[3]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[3]~26 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[3]~26 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[3]~26 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[3]~28 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~105_sumout ),
	.datad(!\D_iw[7]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[3]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[3]~28 .extended_lut = "off";
defparam \R_src1[3]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[3]~28 .shared_arith = "off";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\R_src1[3]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~26_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[4]~0 (
	.dataa(!\E_shift_rot_result[3]~q ),
	.datab(!\E_shift_rot_result[5]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[4]~0 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[4]~0 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[4]~2 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[8]~q ),
	.datad(!\Add0~1_sumout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[4]~2 .extended_lut = "off";
defparam \R_src1[4]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[4]~2 .shared_arith = "off";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\R_src1[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~0_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[1]~0 .extended_lut = "off";
defparam \D_logic_op_raw[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~0 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~0 .lut_mask = 64'hFFFFFFFF6F9F9F6F;
defparam \D_ctrl_alu_force_xor~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~1 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~1 .lut_mask = 64'hFFFFFFFFEFDFDFEF;
defparam \D_ctrl_alu_force_xor~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~3 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~3 .lut_mask = 64'hFFFFFFFFFFFFDF8F;
defparam \D_ctrl_alu_force_xor~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~2 (
	.dataa(!\D_ctrl_alu_force_xor~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~1_combout ),
	.datac(gnd),
	.datad(!\D_ctrl_alu_force_xor~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~2 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~2 .lut_mask = 64'h5533553355335533;
defparam \D_ctrl_alu_force_xor~2 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[1]~0 (
	.dataa(!\D_logic_op_raw[1]~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[1]~0 .extended_lut = "off";
defparam \D_logic_op[1]~0 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[1]~0 .shared_arith = "off";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[0]~1 .extended_lut = "off";
defparam \D_logic_op_raw[0]~1 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[0]~1 (
	.dataa(!\D_ctrl_alu_force_xor~2_combout ),
	.datab(!\D_logic_op_raw[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[0]~1 .extended_lut = "off";
defparam \D_logic_op[0]~1 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[0]~1 .shared_arith = "off";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[4]~0 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[4]~q ),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[4]~0 .extended_lut = "off";
defparam \E_logic_result[4]~0 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~2 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~2 .lut_mask = 64'hFFFFBFFBFFFFBFFB;
defparam \D_ctrl_alu_subtract~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'hFFFFFFD7FFFFFF7D;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'hFFFFDFFDFFFFDFFD;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_sub~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\R_valid~q ),
	.datac(!\D_ctrl_alu_subtract~2_combout ),
	.datad(!\D_ctrl_alu_subtract~1_combout ),
	.datae(!\D_ctrl_alu_subtract~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_sub~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_sub~0 .extended_lut = "off";
defparam \E_alu_sub~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_sub~0 .shared_arith = "off";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cyclonev_lcell_comb \Add2~122 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add2~122_cout ),
	.shareout());
defparam \Add2~122 .extended_lut = "off";
defparam \Add2~122 .lut_mask = 64'h0000000000005555;
defparam \Add2~122 .shared_arith = "off";

cyclonev_lcell_comb \Add2~113 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~q ),
	.datag(gnd),
	.cin(\Add2~122_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~113_sumout ),
	.cout(\Add2~114 ),
	.shareout());
defparam \Add2~113 .extended_lut = "off";
defparam \Add2~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~113 .shared_arith = "off";

cyclonev_lcell_comb \Add2~109 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~q ),
	.datag(gnd),
	.cin(\Add2~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~109_sumout ),
	.cout(\Add2~110 ),
	.shareout());
defparam \Add2~109 .extended_lut = "off";
defparam \Add2~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~109 .shared_arith = "off";

cyclonev_lcell_comb \Add2~101 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~q ),
	.datag(gnd),
	.cin(\Add2~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~101_sumout ),
	.cout(\Add2~102 ),
	.shareout());
defparam \Add2~101 .extended_lut = "off";
defparam \Add2~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~101 .shared_arith = "off";

cyclonev_lcell_comb \Add2~105 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~q ),
	.datag(gnd),
	.cin(\Add2~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~105_sumout ),
	.cout(\Add2~106 ),
	.shareout());
defparam \Add2~105 .extended_lut = "off";
defparam \Add2~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~105 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~q ),
	.datag(gnd),
	.cin(\Add2~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4]~0 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[4]~q ),
	.datad(!\E_logic_result[4]~0_combout ),
	.datae(!\Add2~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4]~0 .extended_lut = "off";
defparam \E_alu_result[4]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~3 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~3 .extended_lut = "off";
defparam \Equal62~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \Equal62~3 .shared_arith = "off";

cyclonev_lcell_comb D_op_rdctl(
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_op_rdctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_op_rdctl.extended_lut = "off";
defparam D_op_rdctl.lut_mask = 64'h7777777777777777;
defparam D_op_rdctl.shared_arith = "off";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal0~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~4 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~4 .extended_lut = "off";
defparam \Equal62~4 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal62~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~5 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~5 .extended_lut = "off";
defparam \Equal62~5 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal62~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_br_cmp~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~3_combout ),
	.datac(!\Equal62~4_combout ),
	.datad(!\Equal62~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br_cmp~0 .extended_lut = "off";
defparam \D_ctrl_br_cmp~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_br_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~7 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~7 .extended_lut = "off";
defparam \Equal0~7 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal0~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~8 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~8 .extended_lut = "off";
defparam \Equal0~8 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal0~8 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_br_cmp~1 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Equal0~8_combout ),
	.datac(!\R_ctrl_br_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br_cmp~1 .extended_lut = "off";
defparam \D_ctrl_br_cmp~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ctrl_br_cmp~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(!\Equal0~1_combout ),
	.datab(!\Equal0~5_combout ),
	.datac(!\Equal0~6_combout ),
	.datad(!\D_ctrl_br_cmp~0_combout ),
	.datae(!\Equal0~7_combout ),
	.dataf(!\D_ctrl_br_cmp~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br_cmp~2 .extended_lut = "off";
defparam \D_ctrl_br_cmp~2 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \D_ctrl_br_cmp~2 .shared_arith = "off";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cyclonev_lcell_comb \E_alu_result~1 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~1 .extended_lut = "off";
defparam \E_alu_result~1 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[5]~0 (
	.dataa(!\R_ctrl_src_imm5_shift_rot~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[5]~0 .extended_lut = "off";
defparam \E_src2[5]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_src2[5]~0 .shared_arith = "off";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[5]~1 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[5]~q ),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[5]~1 .extended_lut = "off";
defparam \E_logic_result[5]~1 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5]~2 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[5]~q ),
	.datad(!\E_logic_result[5]~1_combout ),
	.datae(!\Add2~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5]~2 .extended_lut = "off";
defparam \E_alu_result[5]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[5]~2 .shared_arith = "off";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[9]~2 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[9]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[9]~2 .extended_lut = "off";
defparam \E_logic_result[9]~2 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[9]~2 .shared_arith = "off";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cyclonev_lcell_comb \Add2~77 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~77_sumout ),
	.cout(\Add2~78 ),
	.shareout());
defparam \Add2~77 .extended_lut = "off";
defparam \Add2~77 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~77 .shared_arith = "off";

cyclonev_lcell_comb \Add2~81 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~q ),
	.datag(gnd),
	.cin(\Add2~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~81_sumout ),
	.cout(\Add2~82 ),
	.shareout());
defparam \Add2~81 .extended_lut = "off";
defparam \Add2~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~81 .shared_arith = "off";

cyclonev_lcell_comb \Add2~85 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~q ),
	.datag(gnd),
	.cin(\Add2~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~85_sumout ),
	.cout(\Add2~86 ),
	.shareout());
defparam \Add2~85 .extended_lut = "off";
defparam \Add2~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~85 .shared_arith = "off";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~q ),
	.datag(gnd),
	.cin(\Add2~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~3 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[9]~q ),
	.datad(!\E_logic_result[9]~2_combout ),
	.datae(!\Add2~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~3 .extended_lut = "off";
defparam \E_alu_result[9]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[9]~3 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[8]~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[8]~0 .extended_lut = "off";
defparam \R_src2_hi[8]~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~2 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~2 .extended_lut = "off";
defparam \D_ctrl_logic~2 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \D_ctrl_logic~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_unsigned_lo_imm16~0 (
	.dataa(!\Equal0~1_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\R_src2_use_imm~1_combout ),
	.datad(!\D_ctrl_logic~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_unsigned_lo_imm16~0 .extended_lut = "off";
defparam \D_ctrl_unsigned_lo_imm16~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_unsigned_lo_imm16~0 .shared_arith = "off";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cyclonev_lcell_comb \R_src2_hi~1 (
	.dataa(!\R_ctrl_force_src2_zero~q ),
	.datab(!\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi~1 .extended_lut = "off";
defparam \R_src2_hi~1 .lut_mask = 64'h7777777777777777;
defparam \R_src2_hi~1 .shared_arith = "off";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\R_src2_hi[8]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[24]~3 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[24]~q ),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[24]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[24]~3 .extended_lut = "off";
defparam \E_logic_result[24]~3 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[24]~3 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[7]~10 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[7]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[7]~10 .extended_lut = "off";
defparam \R_src2_hi[7]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[7]~10 .shared_arith = "off";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\R_src2_hi[7]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[6]~9 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[6]~9 .extended_lut = "off";
defparam \R_src2_hi[6]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[6]~9 .shared_arith = "off";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\R_src2_hi[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[5]~8 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[5]~8 .extended_lut = "off";
defparam \R_src2_hi[5]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[5]~8 .shared_arith = "off";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\R_src2_hi[5]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[4]~6 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[10]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[4]~6 .extended_lut = "off";
defparam \R_src2_hi[4]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[4]~6 .shared_arith = "off";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\R_src2_hi[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[3]~7 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[9]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[3]~7 .extended_lut = "off";
defparam \R_src2_hi[3]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[3]~7 .shared_arith = "off";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\R_src2_hi[3]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[2]~11 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[2]~11 .extended_lut = "off";
defparam \R_src2_hi[2]~11 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \R_src2_hi[2]~11 .shared_arith = "off";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\R_src2_hi[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[1]~12 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[1]~12 .extended_lut = "off";
defparam \R_src2_hi[1]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[1]~12 .shared_arith = "off";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\R_src2_hi[1]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[0]~13 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[0]~13 .extended_lut = "off";
defparam \R_src2_hi[0]~13 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[0]~13 .shared_arith = "off";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\R_src2_hi[0]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[5]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cyclonev_lcell_comb \Add2~97 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~97_sumout ),
	.cout(\Add2~98 ),
	.shareout());
defparam \Add2~97 .extended_lut = "off";
defparam \Add2~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~97 .shared_arith = "off";

cyclonev_lcell_comb \Add2~93 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(\Add2~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~93_sumout ),
	.cout(\Add2~94 ),
	.shareout());
defparam \Add2~93 .extended_lut = "off";
defparam \Add2~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~93 .shared_arith = "off";

cyclonev_lcell_comb \Add2~89 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(\Add2~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~89_sumout ),
	.cout(\Add2~90 ),
	.shareout());
defparam \Add2~89 .extended_lut = "off";
defparam \Add2~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~89 .shared_arith = "off";

cyclonev_lcell_comb \Add2~73 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~q ),
	.datag(gnd),
	.cin(\Add2~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~73_sumout ),
	.cout(\Add2~74 ),
	.shareout());
defparam \Add2~73 .extended_lut = "off";
defparam \Add2~73 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~73 .shared_arith = "off";

cyclonev_lcell_comb \Add2~69 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(\Add2~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~69_sumout ),
	.cout(\Add2~70 ),
	.shareout());
defparam \Add2~69 .extended_lut = "off";
defparam \Add2~69 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~69 .shared_arith = "off";

cyclonev_lcell_comb \Add2~65 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~q ),
	.datag(gnd),
	.cin(\Add2~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~65_sumout ),
	.cout(\Add2~66 ),
	.shareout());
defparam \Add2~65 .extended_lut = "off";
defparam \Add2~65 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~65 .shared_arith = "off";

cyclonev_lcell_comb \Add2~61 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(\Add2~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~61_sumout ),
	.cout(\Add2~62 ),
	.shareout());
defparam \Add2~61 .extended_lut = "off";
defparam \Add2~61 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~61 .shared_arith = "off";

cyclonev_lcell_comb \Add2~57 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(\Add2~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~57_sumout ),
	.cout(\Add2~58 ),
	.shareout());
defparam \Add2~57 .extended_lut = "off";
defparam \Add2~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~57 .shared_arith = "off";

cyclonev_lcell_comb \Add2~53 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(\Add2~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~53_sumout ),
	.cout(\Add2~54 ),
	.shareout());
defparam \Add2~53 .extended_lut = "off";
defparam \Add2~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~53 .shared_arith = "off";

cyclonev_lcell_comb \Add2~37 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(\Add2~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~37_sumout ),
	.cout(\Add2~38 ),
	.shareout());
defparam \Add2~37 .extended_lut = "off";
defparam \Add2~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~37 .shared_arith = "off";

cyclonev_lcell_comb \Add2~33 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(\Add2~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout());
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~33 .shared_arith = "off";

cyclonev_lcell_comb \Add2~41 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~q ),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~41_sumout ),
	.cout(\Add2~42 ),
	.shareout());
defparam \Add2~41 .extended_lut = "off";
defparam \Add2~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~41 .shared_arith = "off";

cyclonev_lcell_comb \Add2~45 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~q ),
	.datag(gnd),
	.cin(\Add2~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~45_sumout ),
	.cout(\Add2~46 ),
	.shareout());
defparam \Add2~45 .extended_lut = "off";
defparam \Add2~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~45 .shared_arith = "off";

cyclonev_lcell_comb \Add2~49 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(\Add2~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~49_sumout ),
	.cout(\Add2~50 ),
	.shareout());
defparam \Add2~49 .extended_lut = "off";
defparam \Add2~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~49 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~q ),
	.datag(gnd),
	.cin(\Add2~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24]~4 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[24]~q ),
	.datad(!\E_logic_result[24]~3_combout ),
	.datae(!\Add2~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24]~4 .extended_lut = "off";
defparam \E_alu_result[24]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[24]~4 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[9]~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[9]~2 .extended_lut = "off";
defparam \R_src2_hi[9]~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[9]~2 .shared_arith = "off";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\R_src2_hi[9]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[25]~4 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[25]~q ),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[25]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[25]~4 .extended_lut = "off";
defparam \E_logic_result[25]~4 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[25]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add2~17 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25]~5 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[25]~q ),
	.datad(!\E_logic_result[25]~4_combout ),
	.datae(!\Add2~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25]~5 .extended_lut = "off";
defparam \E_alu_result[25]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[25]~5 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[10]~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[10]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[10]~3 .extended_lut = "off";
defparam \R_src2_hi[10]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[10]~3 .shared_arith = "off";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\R_src2_hi[10]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[26]~5 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[26]~q ),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[26]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[26]~5 .extended_lut = "off";
defparam \E_logic_result[26]~5 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[26]~5 .shared_arith = "off";

cyclonev_lcell_comb \Add2~21 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~21 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26]~6 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[26]~q ),
	.datad(!\E_logic_result[26]~5_combout ),
	.datae(!\Add2~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26]~6 .extended_lut = "off";
defparam \E_alu_result[26]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[26]~6 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[11]~4 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[11]~4 .extended_lut = "off";
defparam \R_src2_hi[11]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[11]~4 .shared_arith = "off";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\R_src2_hi[11]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[27]~6 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[27]~q ),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[27]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[27]~6 .extended_lut = "off";
defparam \E_logic_result[27]~6 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[27]~6 .shared_arith = "off";

cyclonev_lcell_comb \Add2~25 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~q ),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~25 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27]~7 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[27]~q ),
	.datad(!\E_logic_result[27]~6_combout ),
	.datae(!\Add2~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27]~7 .extended_lut = "off";
defparam \E_alu_result[27]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[27]~7 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[12]~5 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[12]~5 .extended_lut = "off";
defparam \R_src2_hi[12]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[12]~5 .shared_arith = "off";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\R_src2_hi[12]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[28]~7 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[28]~q ),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[28]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[28]~7 .extended_lut = "off";
defparam \E_logic_result[28]~7 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[28]~7 .shared_arith = "off";

cyclonev_lcell_comb \Add2~29 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~q ),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout());
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~29 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28]~8 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[28]~q ),
	.datad(!\E_logic_result[28]~7_combout ),
	.datae(!\Add2~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28]~8 .extended_lut = "off";
defparam \E_alu_result[28]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[28]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[20]~8 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[20]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[20]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[20]~8 .extended_lut = "off";
defparam \E_logic_result[20]~8 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[20]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20]~9 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[20]~q ),
	.datad(!\E_logic_result[20]~8_combout ),
	.datae(!\Add2~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20]~9 .extended_lut = "off";
defparam \E_alu_result[20]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[20]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[19]~9 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[19]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[19]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[19]~9 .extended_lut = "off";
defparam \E_logic_result[19]~9 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[19]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19]~10 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[19]~q ),
	.datad(!\E_logic_result[19]~9_combout ),
	.datae(!\Add2~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19]~10 .extended_lut = "off";
defparam \E_alu_result[19]~10 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[19]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[21]~10 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[21]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[21]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[21]~10 .extended_lut = "off";
defparam \E_logic_result[21]~10 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[21]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21]~11 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[21]~q ),
	.datad(!\E_logic_result[21]~10_combout ),
	.datae(!\Add2~41_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21]~11 .extended_lut = "off";
defparam \E_alu_result[21]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[21]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[22]~11 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[22]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[22]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[22]~11 .extended_lut = "off";
defparam \E_logic_result[22]~11 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[22]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22]~12 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[22]~q ),
	.datad(!\E_logic_result[22]~11_combout ),
	.datae(!\Add2~45_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22]~12 .extended_lut = "off";
defparam \E_alu_result[22]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[22]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[23]~12 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[23]~q ),
	.datad(!\E_src1[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[23]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[23]~12 .extended_lut = "off";
defparam \E_logic_result[23]~12 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[23]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23]~13 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[23]~q ),
	.datad(!\E_logic_result[23]~12_combout ),
	.datae(!\Add2~49_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23]~13 .extended_lut = "off";
defparam \E_alu_result[23]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[23]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[18]~13 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[18]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[18]~13 .extended_lut = "off";
defparam \E_logic_result[18]~13 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[18]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18]~14 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[18]~q ),
	.datad(!\E_logic_result[18]~13_combout ),
	.datae(!\Add2~53_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18]~14 .extended_lut = "off";
defparam \E_alu_result[18]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[18]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[17]~14 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[17]~q ),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[17]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[17]~14 .extended_lut = "off";
defparam \E_logic_result[17]~14 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[17]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17]~15 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[17]~q ),
	.datad(!\E_logic_result[17]~14_combout ),
	.datae(!\Add2~57_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17]~15 .extended_lut = "off";
defparam \E_alu_result[17]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[17]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[16]~15 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[16]~q ),
	.datad(!\E_src1[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[16]~15 .extended_lut = "off";
defparam \E_logic_result[16]~15 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[16]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[16]~16 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[16]~q ),
	.datad(!\E_logic_result[16]~15_combout ),
	.datae(!\Add2~61_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16]~16 .extended_lut = "off";
defparam \E_alu_result[16]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[16]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[15]~16 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[15]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[15]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[15]~16 .extended_lut = "off";
defparam \E_logic_result[15]~16 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[15]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15]~17 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[15]~q ),
	.datad(!\E_logic_result[15]~16_combout ),
	.datae(!\Add2~65_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15]~17 .extended_lut = "off";
defparam \E_alu_result[15]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[15]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[14]~17 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[14]~q ),
	.datad(!\E_src1[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[14]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[14]~17 .extended_lut = "off";
defparam \E_logic_result[14]~17 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[14]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14]~18 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[14]~q ),
	.datad(!\E_logic_result[14]~17_combout ),
	.datae(!\Add2~69_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14]~18 .extended_lut = "off";
defparam \E_alu_result[14]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[14]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[13]~18 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[13]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[13]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[13]~18 .extended_lut = "off";
defparam \E_logic_result[13]~18 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[13]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13]~19 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[13]~q ),
	.datad(!\E_logic_result[13]~18_combout ),
	.datae(!\Add2~73_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~19 .extended_lut = "off";
defparam \E_alu_result[13]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[13]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[6]~19 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[6]~q ),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[6]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[6]~19 .extended_lut = "off";
defparam \E_logic_result[6]~19 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[6]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6]~20 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[6]~q ),
	.datad(!\E_logic_result[6]~19_combout ),
	.datae(!\Add2~77_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6]~20 .extended_lut = "off";
defparam \E_alu_result[6]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[6]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[7]~20 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[7]~q ),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[7]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[7]~20 .extended_lut = "off";
defparam \E_logic_result[7]~20 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7]~21 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[7]~q ),
	.datad(!\E_logic_result[7]~20_combout ),
	.datae(!\Add2~81_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7]~21 .extended_lut = "off";
defparam \E_alu_result[7]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[7]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[8]~21 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[8]~q ),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[8]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[8]~21 .extended_lut = "off";
defparam \E_logic_result[8]~21 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[8]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~22 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[8]~q ),
	.datad(!\E_logic_result[8]~21_combout ),
	.datae(!\Add2~85_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~22 .extended_lut = "off";
defparam \E_alu_result[8]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[8]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[12]~22 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[12]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[12]~22 .extended_lut = "off";
defparam \E_logic_result[12]~22 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[12]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~23 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[12]~q ),
	.datad(!\E_logic_result[12]~22_combout ),
	.datae(!\Add2~89_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~23 .extended_lut = "off";
defparam \E_alu_result[12]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[12]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[11]~23 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[11]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[11]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[11]~23 .extended_lut = "off";
defparam \E_logic_result[11]~23 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[11]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~24 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[11]~q ),
	.datad(!\E_logic_result[11]~23_combout ),
	.datae(!\Add2~93_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~24 .extended_lut = "off";
defparam \E_alu_result[11]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[11]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[10]~24 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[10]~q ),
	.datad(!\E_src1[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[10]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[10]~24 .extended_lut = "off";
defparam \E_logic_result[10]~24 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[10]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~25 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[10]~q ),
	.datad(!\E_logic_result[10]~24_combout ),
	.datae(!\Add2~97_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~25 .extended_lut = "off";
defparam \E_alu_result[10]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[10]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[2]~25 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_src2[2]~q ),
	.datac(!\R_logic_op[1]~q ),
	.datad(!\R_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[2]~25 .extended_lut = "off";
defparam \E_logic_result[2]~25 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[2]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2]~26 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\E_shift_rot_result[2]~q ),
	.datac(!\R_ctrl_logic~q ),
	.datad(!\E_logic_result[2]~25_combout ),
	.datae(!\Add2~101_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2]~26 .extended_lut = "off";
defparam \E_alu_result[2]~26 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \E_alu_result[2]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[3]~26 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[3]~q ),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[3]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[3]~26 .extended_lut = "off";
defparam \E_logic_result[3]~26 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[3]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3]~27 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[3]~q ),
	.datad(!\E_logic_result[3]~26_combout ),
	.datae(!\Add2~105_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3]~27 .extended_lut = "off";
defparam \E_alu_result[3]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[3]~27 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_sel_nxt.01~0 (
	.dataa(!\R_ctrl_exception~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt.01~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt.01~0 .extended_lut = "off";
defparam \F_pc_sel_nxt.01~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_pc_sel_nxt.01~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~14 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~14 .extended_lut = "off";
defparam \Equal0~14 .lut_mask = 64'hFFFFFFFFFFBFFFFF;
defparam \Equal0~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~2 .extended_lut = "off";
defparam \Equal62~2 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal62~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~2_combout ),
	.datac(!\Equal0~2_combout ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Equal62~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_invert_arith_src_msb~0 .extended_lut = "off";
defparam \E_invert_arith_src_msb~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \E_invert_arith_src_msb~0 .shared_arith = "off";

cyclonev_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(!\R_valid~q ),
	.datab(!\Equal0~8_combout ),
	.datac(!\Equal0~14_combout ),
	.datad(!\E_invert_arith_src_msb~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_invert_arith_src_msb~1 .extended_lut = "off";
defparam \E_invert_arith_src_msb~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_invert_arith_src_msb~1 .shared_arith = "off";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cyclonev_lcell_comb \R_src2_hi[15]~14 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\R_src2_hi~1_combout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[15]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[15]~14 .extended_lut = "off";
defparam \R_src2_hi[15]~14 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \R_src2_hi[15]~14 .shared_arith = "off";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[14]~15 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_iw[20]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[14]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[14]~15 .extended_lut = "off";
defparam \R_src2_hi[14]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[14]~15 .shared_arith = "off";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\R_src2_hi[14]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[13]~16 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_iw[19]~q ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[13]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[13]~16 .extended_lut = "off";
defparam \R_src2_hi[13]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[13]~16 .shared_arith = "off";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\R_src2_hi[13]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclonev_lcell_comb \Add2~117 (
	.dataa(gnd),
	.datab(!\E_alu_sub~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~117_sumout ),
	.cout(),
	.shareout());
defparam \Add2~117 .extended_lut = "off";
defparam \Add2~117 .lut_mask = 64'h0000000000003333;
defparam \Add2~117 .shared_arith = "off";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[31]~27 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[31]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[31]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[31]~27 .extended_lut = "off";
defparam \E_logic_result[31]~27 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[31]~27 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[30]~28 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[30]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[30]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[30]~28 .extended_lut = "off";
defparam \E_logic_result[30]~28 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[30]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[29]~29 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[29]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[29]~29 .extended_lut = "off";
defparam \E_logic_result[29]~29 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[29]~29 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[1]~30 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[1]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[1]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[1]~30 .extended_lut = "off";
defparam \E_logic_result[1]~30 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[1]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[0]~31 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[0]~31 .extended_lut = "off";
defparam \E_logic_result[0]~31 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[0]~31 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~0 (
	.dataa(!\E_logic_result[2]~25_combout ),
	.datab(!\E_logic_result[3]~26_combout ),
	.datac(!\E_logic_result[18]~13_combout ),
	.datad(!\E_logic_result[0]~31_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~0 .extended_lut = "off";
defparam \Equal127~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal127~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~1 (
	.dataa(!\E_logic_result[31]~27_combout ),
	.datab(!\E_logic_result[30]~28_combout ),
	.datac(!\E_logic_result[29]~29_combout ),
	.datad(!\E_logic_result[1]~30_combout ),
	.datae(!\Equal127~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~1 .extended_lut = "off";
defparam \Equal127~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal127~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~2 (
	.dataa(!\E_logic_result[4]~0_combout ),
	.datab(!\E_logic_result[5]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~2 .extended_lut = "off";
defparam \Equal127~2 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal127~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~3 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[20]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(!\E_src2[19]~q ),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~3 .extended_lut = "off";
defparam \Equal127~3 .lut_mask = 64'h6996966996696996;
defparam \Equal127~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~4 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[6]~q ),
	.datad(!\E_src2[6]~q ),
	.datae(!\E_src1[28]~q ),
	.dataf(!\E_src2[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~4 .extended_lut = "off";
defparam \Equal127~4 .lut_mask = 64'h6996966996696996;
defparam \Equal127~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~5 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[26]~q ),
	.datad(!\E_src2[26]~q ),
	.datae(!\E_src1[27]~q ),
	.dataf(!\E_src2[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~5 .extended_lut = "off";
defparam \Equal127~5 .lut_mask = 64'h6996966996696996;
defparam \Equal127~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~6 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[17]~q ),
	.datad(!\E_src2[17]~q ),
	.datae(!\E_src2[16]~q ),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~6 .extended_lut = "off";
defparam \Equal127~6 .lut_mask = 64'h6996966996696996;
defparam \Equal127~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~7 (
	.dataa(!\E_logic_result[24]~3_combout ),
	.datab(!\E_logic_result[25]~4_combout ),
	.datac(!\Equal127~3_combout ),
	.datad(!\Equal127~4_combout ),
	.datae(!\Equal127~5_combout ),
	.dataf(!\Equal127~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~7 .extended_lut = "off";
defparam \Equal127~7 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal127~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~8 (
	.dataa(!\E_logic_result[10]~24_combout ),
	.datab(!\E_logic_result[9]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~8 .extended_lut = "off";
defparam \Equal127~8 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal127~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~9 (
	.dataa(!\E_logic_result[12]~22_combout ),
	.datab(!\E_logic_result[11]~23_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~9 .extended_lut = "off";
defparam \Equal127~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal127~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~10 (
	.dataa(!\E_logic_result[14]~17_combout ),
	.datab(!\E_logic_result[13]~18_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~10 .extended_lut = "off";
defparam \Equal127~10 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal127~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~11 (
	.dataa(!\E_logic_result[7]~20_combout ),
	.datab(!\E_logic_result[8]~21_combout ),
	.datac(!\E_logic_result[15]~16_combout ),
	.datad(!\E_logic_result[21]~10_combout ),
	.datae(!\E_logic_result[22]~11_combout ),
	.dataf(!\E_logic_result[23]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~11 .extended_lut = "off";
defparam \Equal127~11 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal127~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~12 (
	.dataa(!\Equal127~2_combout ),
	.datab(!\Equal127~7_combout ),
	.datac(!\Equal127~8_combout ),
	.datad(!\Equal127~9_combout ),
	.datae(!\Equal127~10_combout ),
	.dataf(!\Equal127~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~12 .extended_lut = "off";
defparam \Equal127~12 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal127~12 .shared_arith = "off";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \E_cmp_result~0 (
	.dataa(!\Add2~117_sumout ),
	.datab(!\R_compare_op[0]~q ),
	.datac(!\Equal127~1_combout ),
	.datad(!\Equal127~12_combout ),
	.datae(!\R_compare_op[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_cmp_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_cmp_result~0 .extended_lut = "off";
defparam \E_cmp_result~0 .lut_mask = 64'h9669699696696996;
defparam \E_cmp_result~0 .shared_arith = "off";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cyclonev_lcell_comb \Equal62~11 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~11 .extended_lut = "off";
defparam \Equal62~11 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \Equal62~11 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(!\Equal62~11_combout ),
	.datab(!\Equal62~12_combout ),
	.datac(!\Equal62~13_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_uncond_cti_non_br~0 .extended_lut = "off";
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ctrl_uncond_cti_non_br~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~14_combout ),
	.datac(!\Equal62~15_combout ),
	.datad(!\D_ctrl_uncond_cti_non_br~0_combout ),
	.datae(!\D_ctrl_jmp_direct~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_uncond_cti_non_br~1 .extended_lut = "off";
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \D_ctrl_uncond_cti_non_br~1 .shared_arith = "off";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \Equal0~4 .shared_arith = "off";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

cyclonev_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(!\W_cmp_result~q ),
	.datab(!\R_ctrl_br~q ),
	.datac(!\R_ctrl_uncond_cti_non_br~q ),
	.datad(!\R_ctrl_br_uncond~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt~0 .extended_lut = "off";
defparam \F_pc_sel_nxt~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \F_pc_sel_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(!\R_ctrl_exception~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(!\F_pc_sel_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt.10~0 .extended_lut = "off";
defparam \F_pc_sel_nxt.10~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \F_pc_sel_nxt.10~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[17]~1 (
	.dataa(!\Add2~37_sumout ),
	.datab(!\Add0~37_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[17]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[17]~1 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[17]~1 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[17]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[16]~2 (
	.dataa(!\Add2~53_sumout ),
	.datab(!\Add0~53_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[16]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[16]~2 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[16]~2 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[16]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[18]~3 (
	.dataa(!\Add2~33_sumout ),
	.datab(!\Add0~33_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[18]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[18]~3 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[18]~3 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[18]~3 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[19]~4 (
	.dataa(!\Add2~41_sumout ),
	.datab(!\Add0~41_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[19]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[19]~4 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[19]~4 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[19]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[20]~5 (
	.dataa(!\Add2~45_sumout ),
	.datab(!\Add0~45_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[20]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[20]~5 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[20]~5 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[20]~5 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[21]~6 (
	.dataa(!\Add2~49_sumout ),
	.datab(!\Add0~49_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[21]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[21]~6 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[21]~6 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[21]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[22]~7 (
	.dataa(!\Add2~13_sumout ),
	.datab(!\Add0~13_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[22]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[22]~7 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[22]~7 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[22]~7 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[23]~8 (
	.dataa(!\Add2~17_sumout ),
	.datab(!\Add0~17_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[23]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[23]~8 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[23]~8 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[23]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[24]~9 (
	.dataa(!\Add2~21_sumout ),
	.datab(!\Add0~21_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[24]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[24]~9 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[24]~9 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[24]~9 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[26]~10 (
	.dataa(!\Add2~29_sumout ),
	.datab(!\Add0~29_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[26]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[26]~10 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[26]~10 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt[26]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[15]~11 (
	.dataa(!\Add2~57_sumout ),
	.datab(!\Add0~57_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[15]~11 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[15]~11 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[14]~12 (
	.dataa(!\Add2~61_sumout ),
	.datab(!\Add0~61_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[14]~12 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[14]~12 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[14]~12 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[9]~13 (
	.dataa(!\Add2~93_sumout ),
	.datab(!\Add0~93_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[9]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[9]~13 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[9]~13 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt[9]~13 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[11]~14 (
	.dataa(!\Add2~73_sumout ),
	.datab(!\Add0~73_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[11]~14 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[11]~14 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[11]~14 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[13]~15 (
	.dataa(!\Add2~65_sumout ),
	.datab(!\Add0~65_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[13]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[13]~15 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[13]~15 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[13]~15 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[12]~16 (
	.dataa(!\Add2~69_sumout ),
	.datab(!\Add0~69_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[12]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[12]~16 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[12]~16 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[12]~16 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[10]~17 (
	.dataa(!\Add2~89_sumout ),
	.datab(!\Add0~89_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[10]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[10]~17 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[10]~17 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[10]~17 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[0]~18 (
	.dataa(!\Add2~101_sumout ),
	.datab(!\Add0~101_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[0]~18 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[0]~18 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[0]~18 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[1]~19 (
	.dataa(!\Add2~105_sumout ),
	.datab(!\Add0~105_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[1]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[1]~19 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[1]~19 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[1]~19 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[2]~20 (
	.dataa(!\Add2~1_sumout ),
	.datab(!\Add0~1_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[2]~20 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[2]~20 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[2]~20 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt~21 (
	.dataa(!\Add2~5_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt~21 .extended_lut = "off";
defparam \F_pc_no_crst_nxt~21 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt~21 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[4]~22 (
	.dataa(!\Add2~77_sumout ),
	.datab(!\Add0~77_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[4]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[4]~22 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[4]~22 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[4]~22 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[5]~23 (
	.dataa(!\Add2~81_sumout ),
	.datab(!\Add0~81_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[5]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[5]~23 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[5]~23 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[5]~23 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[6]~24 (
	.dataa(!\Add2~85_sumout ),
	.datab(!\Add0~85_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[6]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[6]~24 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[6]~24 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[6]~24 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[7]~25 (
	.dataa(!\Add2~9_sumout ),
	.datab(!\Add0~9_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[7]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[7]~25 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[7]~25 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[7]~25 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[8]~26 (
	.dataa(!\Add2~97_sumout ),
	.datab(!\Add0~97_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[8]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[8]~26 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[8]~26 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[8]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem8~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem8~0 .extended_lut = "off";
defparam \D_ctrl_mem8~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_mem8~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem8~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem8~1 .extended_lut = "off";
defparam \D_ctrl_mem8~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_ctrl_mem8~1 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[23]~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem8~0_combout ),
	.datac(!\D_ctrl_mem16~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[23]~0 .extended_lut = "off";
defparam \E_st_data[23]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \E_st_data[23]~0 .shared_arith = "off";

cyclonev_lcell_comb d_read_nxt(
	.dataa(!d_read1),
	.datab(!WideOr11),
	.datac(!\E_ld_stall~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_read_nxt.extended_lut = "off";
defparam d_read_nxt.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam d_read_nxt.shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!i_read1),
	.datab(!\W_valid~q ),
	.datac(!WideOr12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[25]~0 (
	.dataa(!\Add2~25_sumout ),
	.datab(!\Add0~25_sumout ),
	.datac(!\R_ctrl_exception~q ),
	.datad(!\R_ctrl_break~q ),
	.datae(!\F_pc_sel_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[25]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[25]~0 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[25]~0 .lut_mask = 64'hFAFFFCFFFAFFFCFF;
defparam \F_pc_no_crst_nxt[25]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem16~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem16~1 .extended_lut = "off";
defparam \D_ctrl_mem16~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_mem16~1 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hEFFEEFFEEFFEEFFE;
defparam \E_mem_byte_en~0 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[1]~1 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~1 .extended_lut = "off";
defparam \E_mem_byte_en[1]~1 .lut_mask = 64'hBFFBBFFBBFFBBFFB;
defparam \E_mem_byte_en[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[2]~2 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~2 .extended_lut = "off";
defparam \E_mem_byte_en[2]~2 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \E_mem_byte_en[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~3 .extended_lut = "off";
defparam \E_mem_byte_en[3]~3 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \E_mem_byte_en[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\R_ctrl_break~q ),
	.datac(!hbreak_enabled1),
	.datad(!\Equal62~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~0 .extended_lut = "off";
defparam \hbreak_enabled~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \hbreak_enabled~0 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[24]~1 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(!\D_ctrl_mem16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~1 .extended_lut = "off";
defparam \E_st_data[24]~1 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \E_st_data[24]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[25]~2 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(!\D_ctrl_mem16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~2 .extended_lut = "off";
defparam \E_st_data[25]~2 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \E_st_data[25]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[26]~3 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(!\D_ctrl_mem16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~3 .extended_lut = "off";
defparam \E_st_data[26]~3 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \E_st_data[26]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[27]~4 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(!\D_ctrl_mem16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~4 .extended_lut = "off";
defparam \E_st_data[27]~4 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \E_st_data[27]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[28]~5 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(!\D_ctrl_mem16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~5 .extended_lut = "off";
defparam \E_st_data[28]~5 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \E_st_data[28]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[29]~6 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~6 .extended_lut = "off";
defparam \E_st_data[29]~6 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \E_st_data[29]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[30]~7 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~7 .extended_lut = "off";
defparam \E_st_data[30]~7 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \E_st_data[30]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[31]~8 (
	.dataa(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(!\D_ctrl_mem8~1_combout ),
	.datad(!\D_ctrl_mem16~1_combout ),
	.datae(!\sdram_demo_nios2_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~8 .extended_lut = "off";
defparam \E_st_data[31]~8 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \E_st_data[31]~8 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_nios2_oci (
	readdata_0,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_1,
	readdata_4,
	readdata_3,
	readdata_2,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_5,
	readdata_8,
	readdata_10,
	readdata_9,
	readdata_28,
	readdata_21,
	readdata_29,
	readdata_30,
	readdata_31,
	readdata_17,
	readdata_18,
	readdata_27,
	readdata_7,
	readdata_6,
	readdata_20,
	readdata_19,
	sr_0,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	always0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	rf_source_valid,
	hbreak_enabled,
	jtag_break,
	WideOr1,
	address_nxt,
	r_early_rst,
	oci_ienable_0,
	oci_single_step_mode,
	writedata_nxt,
	debugaccess_nxt,
	byteenable_nxt,
	resetrequest,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_1;
output 	readdata_4;
output 	readdata_3;
output 	readdata_2;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_5;
output 	readdata_8;
output 	readdata_10;
output 	readdata_9;
output 	readdata_28;
output 	readdata_21;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
output 	readdata_17;
output 	readdata_18;
output 	readdata_27;
output 	readdata_7;
output 	readdata_6;
output 	readdata_20;
output 	readdata_19;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	always0;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	rf_source_valid;
input 	hbreak_enabled;
output 	jtag_break;
input 	WideOr1;
input 	[8:0] address_nxt;
input 	r_early_rst;
output 	oci_ienable_0;
output 	oci_single_step_mode;
input 	[31:0] writedata_nxt;
input 	debugaccess_nxt;
input 	[3:0] byteenable_nxt;
output 	resetrequest;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_ready~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \write~0_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \address[4]~q ;
wire \address[3]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_avalon_reg|Equal0~1_combout ;
wire \debugaccess~q ;
wire \the_sdram_demo_nios2_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \byteenable[0]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ;
wire \the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[8]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \writedata[22]~q ;
wire \byteenable[2]~q ;
wire \writedata[23]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \writedata[25]~q ;
wire \writedata[26]~q ;
wire \writedata[4]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \writedata[13]~q ;
wire \writedata[14]~q ;
wire \writedata[15]~q ;
wire \writedata[16]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \writedata[5]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \writedata[10]~q ;
wire \writedata[9]~q ;
wire \writedata[28]~q ;
wire \writedata[21]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \writedata[29]~q ;
wire \writedata[30]~q ;
wire \writedata[31]~q ;
wire \writedata[17]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \writedata[18]~q ;
wire \writedata[27]~q ;
wire \writedata[7]~q ;
wire \writedata[6]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_sdram_demo_nios2_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \address[8]~q ;
wire \address[0]~q ;
wire \readdata~0_combout ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;


sdram_demo_sdram_demo_nios2_cpu_nios2_oci_break the_sdram_demo_nios2_cpu_nios2_oci_break(
	.break_readreg_0(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_24(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_20(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_17(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_5(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_21(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_6(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_9(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[8]~q ),
	.jdo_0(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_25(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_21(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_2(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_19(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_6(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[6]~q ),
	.jdo_23(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_16(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_24(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_22(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_13(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_10(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_nios2_oci_debug the_sdram_demo_nios2_cpu_nios2_oci_debug(
	.r_sync_rst(r_sync_rst),
	.monitor_ready1(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_ready~q ),
	.jtag_break1(jtag_break),
	.jdo_34(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_21(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[20]~q ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_go1(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_go~q ),
	.resetrequest1(resetrequest),
	.jdo_23(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_24(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[24]~q ),
	.resetlatch1(\the_sdram_demo_nios2_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_22(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[22]~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_nios2_ocimem the_sdram_demo_nios2_cpu_nios2_ocimem(
	.MonDReg_1(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[1]~q ),
	.q_a_0(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_22(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_4(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_3(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.MonDReg_16(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[16]~q ),
	.q_a_11(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_16(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_5(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_8(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_28(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_21(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_29(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_17(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_18(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_27(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_7(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.MonDReg_24(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_25(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_22(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_20(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_23(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_17(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_13(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_9(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_28(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_21(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_30(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_7(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[6]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[0]~q ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.take_action_ocimem_a(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_35(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_34(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_17(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.address_3(\address[3]~q ),
	.debugaccess(\debugaccess~q ),
	.MonDReg_2(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[27]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_21(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[20]~q ),
	.MonDReg_3(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_29(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_19(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.MonDReg_4(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.MonDReg_27(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[27]~q ),
	.writedata_22(\writedata[22]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_4(\writedata[4]~q ),
	.jdo_23(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_16(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_11(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[11]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_12(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_14(\writedata[14]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_16(\writedata[16]~q ),
	.MonDReg_5(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[5]~q ),
	.writedata_5(\writedata[5]~q ),
	.MonDReg_8(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_10(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[10]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_21(\writedata[21]~q ),
	.MonDReg_29(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[29]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_31(\writedata[31]~q ),
	.writedata_17(\writedata[17]~q ),
	.MonDReg_18(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[18]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_7(\writedata[7]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.jdo_24(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_22(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_13(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_10(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_nios2_avalon_reg the_sdram_demo_nios2_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.address_3(\address[3]~q ),
	.Equal0(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.debugaccess(\debugaccess~q ),
	.take_action_ocireg(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_ienable_0(oci_ienable_0),
	.oci_single_step_mode1(oci_single_step_mode),
	.monitor_error(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_error~q ),
	.oci_reg_readdata_0(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ),
	.oci_ienable_8(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[8]~q ),
	.oci_reg_readdata(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.writedata_3(\writedata[3]~q ),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_debug_slave_wrapper the_sdram_demo_nios2_cpu_debug_slave_wrapper(
	.break_readreg_0(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[1]~q ),
	.break_readreg_2(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_24(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_22(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[22]~q ),
	.break_readreg_20(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_23(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[23]~q ),
	.break_readreg_17(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_13(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_9(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_28(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_21(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_30(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_7(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[6]~q ),
	.break_readreg_5(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_21(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_6(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_9(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_sdram_demo_nios2_cpu_nios2_oci_break|break_readreg[8]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.MonDReg_0(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[0]~q ),
	.monitor_ready(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_0(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.take_action_ocimem_a(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_35(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[3]~q ),
	.hbreak_enabled(hbreak_enabled),
	.jdo_34(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_17(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[25]~q ),
	.MonDReg_2(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_21(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[20]~q ),
	.MonDReg_3(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[33]~q ),
	.monitor_error(\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[18]~q ),
	.MonDReg_4(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_27(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[27]~q ),
	.jdo_23(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_16(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_11(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_8(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_10(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_29(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_18(\the_sdram_demo_nios2_cpu_nios2_ocimem|MonDReg[18]~q ),
	.jdo_24(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[7]~q ),
	.resetlatch(\the_sdram_demo_nios2_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_22(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_13(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_10(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_sdram_demo_nios2_cpu_debug_slave_wrapper|the_sdram_demo_nios2_cpu_debug_slave_sysclk|jdo[9]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!always0),
	.datab(!saved_grant_0),
	.datac(!waitrequest),
	.datad(!mem_used_1),
	.datae(!WideOr1),
	.dataf(!\write~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFF3FFFFF7F7FFFFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!\read~q ),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \read~0 .shared_arith = "off";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

cyclonev_lcell_comb \readdata~0 (
	.dataa(!\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_ready~q ),
	.datab(!\address[0]~q ),
	.datac(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~0 .extended_lut = "off";
defparam \readdata~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \readdata~1 (
	.dataa(!\address[0]~q ),
	.datab(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datac(!oci_single_step_mode),
	.datad(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~1 .extended_lut = "off";
defparam \readdata~1 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!\address[0]~q ),
	.datab(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datac(!\the_sdram_demo_nios2_cpu_nios2_avalon_reg|oci_ienable[8]~q ),
	.datad(!\the_sdram_demo_nios2_cpu_nios2_oci_debug|monitor_go~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~2 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_debug_slave_wrapper (
	break_readreg_0,
	break_readreg_1,
	MonDReg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	break_readreg_26,
	MonDReg_26,
	MonDReg_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_23,
	break_readreg_17,
	MonDReg_17,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_9,
	MonDReg_28,
	MonDReg_21,
	MonDReg_30,
	MonDReg_31,
	MonDReg_7,
	MonDReg_6,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_21,
	break_readreg_18,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_9,
	break_readreg_8,
	sr_0,
	ir_out_0,
	ir_out_1,
	MonDReg_0,
	monitor_ready,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	take_action_ocimem_a,
	jdo_35,
	take_action_ocimem_b,
	jdo_3,
	hbreak_enabled,
	jdo_34,
	jdo_17,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_25,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	MonDReg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	monitor_error,
	jdo_19,
	jdo_18,
	MonDReg_4,
	jdo_6,
	MonDReg_27,
	jdo_23,
	jdo_16,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_8,
	MonDReg_10,
	MonDReg_29,
	MonDReg_18,
	jdo_24,
	jdo_7,
	resetlatch,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_10,
	jdo_9,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	break_readreg_1;
input 	MonDReg_1;
input 	break_readreg_2;
input 	break_readreg_3;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	MonDReg_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_23;
input 	break_readreg_17;
input 	MonDReg_17;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_9;
input 	MonDReg_28;
input 	MonDReg_21;
input 	MonDReg_30;
input 	MonDReg_31;
input 	MonDReg_7;
input 	MonDReg_6;
input 	break_readreg_5;
input 	break_readreg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	break_readreg_31;
input 	break_readreg_21;
input 	break_readreg_18;
input 	break_readreg_6;
input 	break_readreg_22;
input 	break_readreg_15;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_9;
input 	break_readreg_8;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	MonDReg_0;
input 	monitor_ready;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	take_action_ocimem_a;
output 	jdo_35;
output 	take_action_ocimem_b;
output 	jdo_3;
input 	hbreak_enabled;
output 	jdo_34;
output 	jdo_17;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	jdo_25;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_21;
output 	jdo_20;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
input 	monitor_error;
output 	jdo_19;
output 	jdo_18;
input 	MonDReg_4;
output 	jdo_6;
input 	MonDReg_27;
output 	jdo_23;
output 	jdo_16;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_8;
input 	MonDReg_10;
input 	MonDReg_29;
input 	MonDReg_18;
output 	jdo_24;
output 	jdo_7;
input 	resetlatch;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_11;
output 	jdo_13;
output 	jdo_12;
output 	jdo_10;
output 	jdo_9;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[1]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[2]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[3]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[4]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[17]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[25]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[5]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[26]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[28]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[27]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[21]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[20]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[18]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[6]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[29]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[30]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[32]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[22]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[19]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[23]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[16]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[24]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[8]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[14]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[11]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[13]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[12]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[10]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[9]~q ;
wire \sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_uir~combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[36]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[37]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[35]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[34]~q ;
wire \sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[31]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[33]~q ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[7]~q ;
wire \sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_sdram_demo_nios2_cpu_debug_slave_tck|sr[15]~q ;


sdram_demo_sdram_demo_nios2_cpu_debug_slave_sysclk the_sdram_demo_nios2_cpu_debug_slave_sysclk(
	.sr_1(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[2]~q ),
	.sr_3(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[3]~q ),
	.sr_4(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[4]~q ),
	.sr_17(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[5]~q ),
	.sr_26(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[27]~q ),
	.sr_21(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[18]~q ),
	.sr_6(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[6]~q ),
	.sr_29(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[29]~q ),
	.sr_30(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[32]~q ),
	.sr_22(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[22]~q ),
	.sr_19(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[19]~q ),
	.sr_23(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[23]~q ),
	.sr_16(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[16]~q ),
	.sr_24(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[24]~q ),
	.sr_8(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[8]~q ),
	.sr_14(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[14]~q ),
	.sr_11(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[11]~q ),
	.sr_13(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[12]~q ),
	.sr_10(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[9]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.jdo_3(jdo_3),
	.jdo_34(jdo_34),
	.jdo_17(jdo_17),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[37]~q ),
	.sr_35(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[35]~q ),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.sr_34(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[34]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_6(jdo_6),
	.sr_31(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[33]~q ),
	.jdo_23(jdo_23),
	.jdo_16(jdo_16),
	.jdo_24(jdo_24),
	.sr_7(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.virtual_state_udr(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_22(jdo_22),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_8(jdo_8),
	.jdo_11(jdo_11),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_15(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[15]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

sdram_demo_sdram_demo_nios2_cpu_debug_slave_tck the_sdram_demo_nios2_cpu_debug_slave_tck(
	.sr_1(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.sr_3(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.sr_4(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.sr_17(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_26(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[27]~q ),
	.sr_21(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.sr_29(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[29]~q ),
	.break_readreg_27(break_readreg_27),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.sr_30(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[32]~q ),
	.MonDReg_22(MonDReg_22),
	.sr_22(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[19]~q ),
	.MonDReg_23(MonDReg_23),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_15(MonDReg_15),
	.MonDReg_9(MonDReg_9),
	.MonDReg_28(MonDReg_28),
	.MonDReg_21(MonDReg_21),
	.MonDReg_30(MonDReg_30),
	.MonDReg_31(MonDReg_31),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.break_readreg_29(break_readreg_29),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.sr_23(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.break_readreg_18(break_readreg_18),
	.sr_16(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[16]~q ),
	.sr_24(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[24]~q ),
	.sr_8(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.break_readreg_22(break_readreg_22),
	.break_readreg_15(break_readreg_15),
	.sr_14(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[14]~q ),
	.sr_11(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[11]~q ),
	.sr_13(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[12]~q ),
	.sr_10(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_23(break_readreg_23),
	.break_readreg_7(break_readreg_7),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_10(break_readreg_10),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_9(break_readreg_9),
	.break_readreg_8(break_readreg_8),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.monitor_ready(monitor_ready),
	.hbreak_enabled(hbreak_enabled),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[37]~q ),
	.sr_35(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[35]~q ),
	.sr_34(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[34]~q ),
	.MonDReg_3(MonDReg_3),
	.virtual_state_cdr(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.monitor_error(monitor_error),
	.MonDReg_4(MonDReg_4),
	.MonDReg_27(MonDReg_27),
	.sr_31(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[33]~q ),
	.MonDReg_11(MonDReg_11),
	.MonDReg_12(MonDReg_12),
	.MonDReg_5(MonDReg_5),
	.MonDReg_8(MonDReg_8),
	.MonDReg_10(MonDReg_10),
	.MonDReg_29(MonDReg_29),
	.MonDReg_18(MonDReg_18),
	.sr_7(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[7]~q ),
	.resetlatch(resetlatch),
	.sr_15(\the_sdram_demo_nios2_cpu_debug_slave_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

sdram_demo_sld_virtual_jtag_basic_1 sdram_demo_nios2_cpu_debug_slave_phy(
	.virtual_state_sdr(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\sdram_demo_nios2_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

endmodule

module sdram_demo_sdram_demo_nios2_cpu_debug_slave_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_4,
	sr_17,
	sr_25,
	sr_5,
	sr_26,
	sr_28,
	sr_27,
	sr_21,
	sr_20,
	sr_18,
	sr_6,
	sr_29,
	sr_30,
	sr_32,
	sr_22,
	sr_19,
	sr_23,
	sr_16,
	sr_24,
	sr_8,
	sr_14,
	sr_11,
	sr_13,
	sr_12,
	sr_10,
	sr_9,
	sr_0,
	virtual_state_uir,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe1,
	take_action_ocimem_a1,
	jdo_35,
	take_action_ocimem_b1,
	jdo_3,
	jdo_34,
	jdo_17,
	take_action_ocimem_a2,
	take_action_ocimem_a3,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	sr_35,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	sr_34,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	jdo_6,
	sr_31,
	sr_33,
	jdo_23,
	jdo_16,
	jdo_24,
	sr_7,
	jdo_7,
	virtual_state_udr,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_10,
	jdo_9,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_4;
input 	sr_17;
input 	sr_25;
input 	sr_5;
input 	sr_26;
input 	sr_28;
input 	sr_27;
input 	sr_21;
input 	sr_20;
input 	sr_18;
input 	sr_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_22;
input 	sr_19;
input 	sr_23;
input 	sr_16;
input 	sr_24;
input 	sr_8;
input 	sr_14;
input 	sr_11;
input 	sr_13;
input 	sr_12;
input 	sr_10;
input 	sr_9;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	take_action_ocimem_a1;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	jdo_3;
output 	jdo_34;
output 	jdo_17;
output 	take_action_ocimem_a2;
output 	take_action_ocimem_a3;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
input 	sr_35;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_21;
output 	jdo_20;
input 	sr_34;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_19;
output 	jdo_18;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
output 	jdo_23;
output 	jdo_16;
output 	jdo_24;
input 	sr_7;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_11;
output 	jdo_13;
output 	jdo_12;
output 	jdo_10;
output 	jdo_9;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


sdram_demo_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

sdram_demo_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cyclonev_lcell_comb take_action_ocimem_b(
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_35),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_b1),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_b.extended_lut = "off";
defparam take_action_ocimem_b.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam take_action_ocimem_b.shared_arith = "off";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(!jdo_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!take_action_ocimem_a2),
	.datab(!jdo_34),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module sdram_demo_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module sdram_demo_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_debug_slave_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	sr_4,
	break_readreg_2,
	sr_17,
	sr_25,
	sr_5,
	break_readreg_3,
	sr_26,
	sr_28,
	sr_27,
	sr_21,
	sr_20,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	sr_29,
	break_readreg_27,
	break_readreg_26,
	MonDReg_26,
	sr_30,
	sr_32,
	MonDReg_22,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	MonDReg_23,
	break_readreg_17,
	MonDReg_17,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_9,
	MonDReg_28,
	MonDReg_21,
	MonDReg_30,
	MonDReg_31,
	MonDReg_7,
	MonDReg_6,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	sr_23,
	break_readreg_21,
	break_readreg_18,
	sr_16,
	sr_24,
	sr_8,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	sr_14,
	sr_11,
	sr_13,
	sr_12,
	sr_10,
	sr_9,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_9,
	break_readreg_8,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	MonDReg_0,
	virtual_state_uir,
	monitor_ready,
	hbreak_enabled,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_35,
	sr_34,
	MonDReg_3,
	virtual_state_cdr,
	monitor_error,
	MonDReg_4,
	MonDReg_27,
	sr_31,
	sr_33,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_8,
	MonDReg_10,
	MonDReg_29,
	MonDReg_18,
	sr_7,
	resetlatch,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
output 	sr_4;
input 	break_readreg_2;
output 	sr_17;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
output 	sr_26;
output 	sr_28;
output 	sr_27;
output 	sr_21;
output 	sr_20;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
output 	sr_29;
input 	break_readreg_27;
input 	break_readreg_26;
input 	MonDReg_26;
output 	sr_30;
output 	sr_32;
input 	MonDReg_22;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
input 	MonDReg_23;
input 	break_readreg_17;
input 	MonDReg_17;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_9;
input 	MonDReg_28;
input 	MonDReg_21;
input 	MonDReg_30;
input 	MonDReg_31;
input 	MonDReg_7;
input 	MonDReg_6;
input 	break_readreg_5;
input 	break_readreg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	break_readreg_31;
output 	sr_23;
input 	break_readreg_21;
input 	break_readreg_18;
output 	sr_16;
output 	sr_24;
output 	sr_8;
input 	break_readreg_6;
input 	break_readreg_22;
input 	break_readreg_15;
output 	sr_14;
output 	sr_11;
output 	sr_13;
output 	sr_12;
output 	sr_10;
output 	sr_9;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_9;
input 	break_readreg_8;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	MonDReg_0;
input 	virtual_state_uir;
input 	monitor_ready;
input 	hbreak_enabled;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_35;
output 	sr_34;
input 	MonDReg_3;
input 	virtual_state_cdr;
input 	monitor_error;
input 	MonDReg_4;
input 	MonDReg_27;
output 	sr_31;
output 	sr_33;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_8;
input 	MonDReg_10;
input 	MonDReg_29;
input 	MonDReg_18;
output 	sr_7;
input 	resetlatch;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[14]~9_combout ;
wire \sr[14]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~13_combout ;
wire \sr~20_combout ;
wire \sr[21]~21_combout ;
wire \sr[21]~19_combout ;
wire \sr~22_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~37_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \sr~14_combout ;
wire \sr[37]~15_combout ;
wire \sr~16_combout ;
wire \Mux37~0_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr[21]~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~38_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr[21]~55_combout ;
wire \DRsize.010~q ;
wire \sr~48_combout ;
wire \sr~49_combout ;


sdram_demo_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

sdram_demo_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[21]~21_combout ),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~15_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~15_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[21]~19_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[14]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[14]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[14]~9 .extended_lut = "off";
defparam \sr[14]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[14]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[14]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[14]~10 .extended_lut = "off";
defparam \sr[14]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[14]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~13 .shared_arith = "off";

cyclonev_lcell_comb \sr~20 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~20 .extended_lut = "off";
defparam \sr~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~20 .shared_arith = "off";

cyclonev_lcell_comb \sr[21]~21 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[21]~21 .extended_lut = "off";
defparam \sr[21]~21 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \sr[21]~19 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[21]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[21]~19 .extended_lut = "off";
defparam \sr[21]~19 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[21]~19 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_19),
	.datad(!break_readreg_17),
	.datae(!MonDReg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_5),
	.datad(!sr_7),
	.datae(!break_readreg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_30),
	.datad(!MonDReg_28),
	.datae(!break_readreg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~32 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_31),
	.datad(!MonDReg_29),
	.datae(!break_readreg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~32 .extended_lut = "off";
defparam \sr~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_33),
	.datad(!MonDReg_31),
	.datae(!break_readreg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_21),
	.datad(!sr_23),
	.datae(!break_readreg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_20),
	.datad(!MonDReg_18),
	.datae(!break_readreg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_22),
	.datad(!sr_24),
	.datae(!break_readreg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_17),
	.datad(!MonDReg_15),
	.datae(!break_readreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_25),
	.datad(!MonDReg_23),
	.datae(!break_readreg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_7),
	.datad(!sr_9),
	.datae(!break_readreg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~50 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~51 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~54 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \sr~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~14 .extended_lut = "off";
defparam \sr~14 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~14 .shared_arith = "off";

cyclonev_lcell_comb \sr[37]~15 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[37]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[37]~15 .extended_lut = "off";
defparam \sr[37]~15 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[37]~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_2),
	.datad(!irf_reg_1_2),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~17 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~17 .extended_lut = "off";
defparam \sr~17 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~17 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr[21]~33 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[21]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[21]~33 .extended_lut = "off";
defparam \sr[21]~33 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[21]~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'h2727272727272727;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~35 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~35 .extended_lut = "off";
defparam \sr~35 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~36 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[21]~33_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~34_combout ),
	.dataf(!\sr~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~36 .extended_lut = "off";
defparam \sr~36 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_6),
	.datac(!break_readreg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h2727272727272727;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_2),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr[21]~55 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[21]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[21]~55 .extended_lut = "off";
defparam \sr[21]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[21]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[21]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_2),
	.datac(!irf_reg_1_2),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~48_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~49 .shared_arith = "off";

endmodule

module sdram_demo_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module sdram_demo_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module sdram_demo_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	writedata_0,
	address_0,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	address_3,
	Equal0,
	debugaccess,
	take_action_ocireg,
	oci_ienable_0,
	oci_single_step_mode1,
	monitor_error,
	oci_reg_readdata_0,
	oci_ienable_8,
	oci_reg_readdata,
	writedata_3,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
input 	writedata_0;
input 	address_0;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	address_3;
output 	Equal0;
input 	debugaccess;
output 	take_action_ocireg;
output 	oci_ienable_0;
output 	oci_single_step_mode1;
input 	monitor_error;
output 	oci_reg_readdata_0;
output 	oci_ienable_8;
output 	oci_reg_readdata;
input 	writedata_3;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \oci_ienable[0]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_single_step_mode~0_combout ;


cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_2),
	.datab(!address_1),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!write),
	.datab(!address_0),
	.datac(!Equal0),
	.datad(!debugaccess),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(\oci_ienable[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata[0]~0 (
	.dataa(!address_0),
	.datab(!Equal0),
	.datac(!oci_ienable_0),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata[0]~0 .extended_lut = "off";
defparam \oci_reg_readdata[0]~0 .lut_mask = 64'hB1FFB1FFB1FFB1FF;
defparam \oci_reg_readdata[0]~0 .shared_arith = "off";

dffeas \oci_ienable[8] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_8),
	.prn(vcc));
defparam \oci_ienable[8] .is_wysiwyg = "true";
defparam \oci_ienable[8] .power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata~1 (
	.dataa(!address_0),
	.datab(!Equal0),
	.datac(!oci_ienable_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~1 .extended_lut = "off";
defparam \oci_reg_readdata~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \oci_reg_readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(!address_4),
	.dataf(!address_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[0]~0 (
	.dataa(!writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[0]~0 .extended_lut = "off";
defparam \oci_ienable[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(!write),
	.datab(!address_0),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(!debugaccess),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_oci_intr_mask_reg~0 .extended_lut = "off";
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam \take_action_oci_intr_mask_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!take_action_ocireg),
	.datab(!oci_single_step_mode1),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h2727272727272727;
defparam \oci_single_step_mode~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_16,
	break_readreg_24,
	break_readreg_4,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_20,
	break_readreg_19,
	break_readreg_17,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_21,
	break_readreg_18,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_9,
	break_readreg_8,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_3,
	jdo_17,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_19,
	jdo_18,
	jdo_6,
	jdo_23,
	jdo_16,
	jdo_24,
	jdo_7,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_3;
output 	break_readreg_16;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_17;
output 	break_readreg_5;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_6;
output 	break_readreg_22;
output 	break_readreg_15;
output 	break_readreg_23;
output 	break_readreg_7;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_10;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_9;
output 	break_readreg_8;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_17;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_21;
input 	jdo_20;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_19;
input 	jdo_18;
input 	jdo_6;
input 	jdo_23;
input 	jdo_16;
input 	jdo_24;
input 	jdo_7;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_11;
input 	jdo_13;
input 	jdo_12;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[23]~0_combout ;
wire \break_readreg[23]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[23]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[23]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

cyclonev_lcell_comb \break_readreg[23]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[23]~0 .extended_lut = "off";
defparam \break_readreg[23]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[23]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[23]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[23]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[23]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[23]~1 .extended_lut = "off";
defparam \break_readreg[23]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[23]~1 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_nios2_oci_debug (
	r_sync_rst,
	monitor_ready1,
	jtag_break1,
	jdo_34,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_25,
	writedata_0,
	take_action_ocireg,
	jdo_21,
	jdo_20,
	writedata_1,
	monitor_error1,
	jdo_19,
	jdo_18,
	monitor_go1,
	resetrequest1,
	jdo_23,
	jdo_24,
	resetlatch1,
	jdo_22,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	monitor_ready1;
output 	jtag_break1;
input 	jdo_34;
input 	take_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_25;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_21;
input 	jdo_20;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_go1;
output 	resetrequest1;
input 	jdo_23;
input 	jdo_24;
output 	resetlatch1;
input 	jdo_22;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \monitor_ready~0_combout ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


sdram_demo_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetrequest(
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(resetrequest1),
	.prn(vcc));
defparam resetrequest.is_wysiwyg = "true";
defparam resetrequest.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!monitor_ready1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_25),
	.datad(!writedata_0),
	.datae(!take_action_ocireg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!\break_on_reset~q ),
	.datab(!jdo_19),
	.datac(!jdo_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_25),
	.datac(!take_action_ocireg),
	.datad(!writedata_1),
	.datae(!monitor_error1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_34),
	.datac(!monitor_go1),
	.datad(!jdo_23),
	.datae(!state_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \monitor_go~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

endmodule

module sdram_demo_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_nios2_ocimem (
	MonDReg_1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_4,
	q_a_3,
	MonDReg_16,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_5,
	q_a_8,
	q_a_10,
	q_a_9,
	q_a_28,
	q_a_21,
	q_a_29,
	q_a_30,
	q_a_31,
	q_a_17,
	q_a_18,
	q_a_27,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	MonDReg_24,
	MonDReg_25,
	MonDReg_26,
	MonDReg_22,
	MonDReg_20,
	MonDReg_19,
	MonDReg_23,
	MonDReg_17,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_9,
	MonDReg_28,
	MonDReg_21,
	MonDReg_30,
	MonDReg_31,
	MonDReg_7,
	MonDReg_6,
	waitrequest1,
	MonDReg_0,
	write,
	address_8,
	read,
	take_action_ocimem_a,
	jdo_35,
	take_action_ocimem_b,
	jdo_3,
	jdo_34,
	jdo_17,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_25,
	writedata_0,
	address_0,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	address_3,
	debugaccess,
	MonDReg_2,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	r_early_rst,
	byteenable_0,
	jdo_21,
	jdo_20,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	writedata_3,
	MonDReg_4,
	jdo_6,
	writedata_2,
	MonDReg_27,
	writedata_22,
	byteenable_2,
	writedata_23,
	writedata_24,
	byteenable_3,
	writedata_25,
	writedata_26,
	writedata_4,
	jdo_23,
	jdo_16,
	MonDReg_11,
	writedata_11,
	byteenable_1,
	MonDReg_12,
	writedata_12,
	writedata_13,
	writedata_14,
	writedata_15,
	writedata_16,
	MonDReg_5,
	writedata_5,
	MonDReg_8,
	writedata_8,
	MonDReg_10,
	writedata_10,
	writedata_9,
	writedata_28,
	writedata_21,
	MonDReg_29,
	writedata_29,
	writedata_30,
	writedata_31,
	writedata_17,
	MonDReg_18,
	writedata_18,
	writedata_27,
	writedata_7,
	writedata_6,
	writedata_20,
	writedata_19,
	jdo_24,
	jdo_7,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_4;
output 	q_a_3;
output 	MonDReg_16;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_5;
output 	q_a_8;
output 	q_a_10;
output 	q_a_9;
output 	q_a_28;
output 	q_a_21;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	q_a_17;
output 	q_a_18;
output 	q_a_27;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_19;
output 	MonDReg_24;
output 	MonDReg_25;
output 	MonDReg_26;
output 	MonDReg_22;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_23;
output 	MonDReg_17;
output 	MonDReg_13;
output 	MonDReg_14;
output 	MonDReg_15;
output 	MonDReg_9;
output 	MonDReg_28;
output 	MonDReg_21;
output 	MonDReg_30;
output 	MonDReg_31;
output 	MonDReg_7;
output 	MonDReg_6;
output 	waitrequest1;
output 	MonDReg_0;
input 	write;
input 	address_8;
input 	read;
input 	take_action_ocimem_a;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	jdo_3;
input 	jdo_34;
input 	jdo_17;
input 	take_action_ocimem_a1;
input 	take_action_ocimem_a2;
input 	jdo_25;
input 	writedata_0;
input 	address_0;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	address_3;
input 	debugaccess;
output 	MonDReg_2;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	r_early_rst;
input 	byteenable_0;
input 	jdo_21;
input 	jdo_20;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
output 	MonDReg_4;
input 	jdo_6;
input 	writedata_2;
output 	MonDReg_27;
input 	writedata_22;
input 	byteenable_2;
input 	writedata_23;
input 	writedata_24;
input 	byteenable_3;
input 	writedata_25;
input 	writedata_26;
input 	writedata_4;
input 	jdo_23;
input 	jdo_16;
output 	MonDReg_11;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_12;
input 	writedata_12;
input 	writedata_13;
input 	writedata_14;
input 	writedata_15;
input 	writedata_16;
output 	MonDReg_5;
input 	writedata_5;
output 	MonDReg_8;
input 	writedata_8;
output 	MonDReg_10;
input 	writedata_10;
input 	writedata_9;
input 	writedata_28;
input 	writedata_21;
output 	MonDReg_29;
input 	writedata_29;
input 	writedata_30;
input 	writedata_31;
input 	writedata_17;
output 	MonDReg_18;
input 	writedata_18;
input 	writedata_27;
input 	writedata_7;
input 	writedata_6;
input 	writedata_20;
input 	writedata_19;
input 	jdo_24;
input 	jdo_7;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_11;
input 	jdo_13;
input 	jdo_12;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[22]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[23]~4_combout ;
wire \ociram_wr_data[24]~5_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~6_combout ;
wire \ociram_wr_data[26]~7_combout ;
wire \ociram_wr_data[4]~8_combout ;
wire \ociram_wr_data[3]~9_combout ;
wire \ociram_wr_data[11]~10_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[12]~11_combout ;
wire \ociram_wr_data[13]~12_combout ;
wire \ociram_wr_data[14]~13_combout ;
wire \ociram_wr_data[15]~14_combout ;
wire \ociram_wr_data[16]~15_combout ;
wire \ociram_wr_data[5]~16_combout ;
wire \ociram_wr_data[8]~17_combout ;
wire \ociram_wr_data[10]~18_combout ;
wire \ociram_wr_data[9]~19_combout ;
wire \ociram_wr_data[28]~20_combout ;
wire \ociram_wr_data[21]~21_combout ;
wire \ociram_wr_data[29]~22_combout ;
wire \ociram_wr_data[30]~23_combout ;
wire \ociram_wr_data[31]~24_combout ;
wire \ociram_wr_data[17]~25_combout ;
wire \ociram_wr_data[18]~26_combout ;
wire \ociram_wr_data[27]~27_combout ;
wire \ociram_wr_data[7]~28_combout ;
wire \ociram_wr_data[6]~29_combout ;
wire \ociram_wr_data[20]~30_combout ;
wire \ociram_wr_data[19]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~5_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~10 ;
wire \Add0~21_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~34 ;
wire \Add0~17_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[9]~3_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~2_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~0_combout ;
wire \MonDReg~1_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg[27]~16_combout ;
wire \MonDReg[27]~7_combout ;
wire \MonDReg[27]~8_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~11_combout ;
wire \MonDReg[8]~12_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~15_combout ;


sdram_demo_sdram_demo_nios2_cpu_ociram_sp_ram_module sdram_demo_nios2_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_4(q_a_4),
	.q_a_3(q_a_3),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_16(q_a_16),
	.q_a_5(q_a_5),
	.q_a_8(q_a_8),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_28(q_a_28),
	.q_a_21(q_a_21),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.q_a_17(q_a_17),
	.q_a_18(q_a_18),
	.q_a_27(q_a_27),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~4_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~5_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~6_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~7_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~8_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~9_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~10_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~11_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~12_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~13_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~14_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~15_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~16_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~17_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~18_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~19_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~20_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~21_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~22_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~23_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~24_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~25_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~26_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~27_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~28_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~29_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~30_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!write),
	.datab(!address_8),
	.datac(!\jtag_ram_access~q ),
	.datad(!debugaccess),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!address_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[5]~q ),
	.datac(!address_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[6]~q ),
	.datac(!address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[7]~q ),
	.datac(!address_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[8]~q ),
	.datac(!address_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[9]~q ),
	.datac(!address_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_1),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\Add0~1_sumout ),
	.datad(!\jtag_ram_wr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~3 .extended_lut = "off";
defparam \ociram_wr_data[22]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~1 .extended_lut = "off";
defparam \ociram_byteenable[2]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~4 .extended_lut = "off";
defparam \ociram_wr_data[23]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~5 .extended_lut = "off";
defparam \ociram_wr_data[24]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~2 .extended_lut = "off";
defparam \ociram_byteenable[3]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~6 .extended_lut = "off";
defparam \ociram_wr_data[25]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~7 .extended_lut = "off";
defparam \ociram_wr_data[26]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~8 .extended_lut = "off";
defparam \ociram_wr_data[4]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_3),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~9 .extended_lut = "off";
defparam \ociram_wr_data[3]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[3]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~10 .extended_lut = "off";
defparam \ociram_wr_data[11]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~3 .extended_lut = "off";
defparam \ociram_byteenable[1]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~11 .extended_lut = "off";
defparam \ociram_wr_data[12]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~12 .extended_lut = "off";
defparam \ociram_wr_data[13]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~13 .extended_lut = "off";
defparam \ociram_wr_data[14]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~14 .extended_lut = "off";
defparam \ociram_wr_data[15]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_16),
	.datac(!writedata_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~15 .extended_lut = "off";
defparam \ociram_wr_data[16]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~16 .extended_lut = "off";
defparam \ociram_wr_data[5]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~17 .extended_lut = "off";
defparam \ociram_wr_data[8]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~18 .extended_lut = "off";
defparam \ociram_wr_data[10]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~19 .extended_lut = "off";
defparam \ociram_wr_data[9]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~20 .extended_lut = "off";
defparam \ociram_wr_data[28]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~21 .extended_lut = "off";
defparam \ociram_wr_data[21]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~22 .extended_lut = "off";
defparam \ociram_wr_data[29]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~23 .extended_lut = "off";
defparam \ociram_wr_data[30]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~24 .extended_lut = "off";
defparam \ociram_wr_data[31]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~25 .extended_lut = "off";
defparam \ociram_wr_data[17]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~26 .extended_lut = "off";
defparam \ociram_wr_data[18]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~27 .extended_lut = "off";
defparam \ociram_wr_data[27]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~28 .extended_lut = "off";
defparam \ociram_wr_data[7]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~29 .extended_lut = "off";
defparam \ociram_wr_data[6]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~30 .extended_lut = "off";
defparam \ociram_wr_data[20]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~31 .extended_lut = "off";
defparam \ociram_wr_data[19]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~31 .shared_arith = "off";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(q_a_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(q_a_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(q_a_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(q_a_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(q_a_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(q_a_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[9]~3_combout ),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(\MonDReg[27]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[27]~8_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[27]~8_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_34),
	.datac(!jdo_17),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_b),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[9]~3 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[9]~3 .extended_lut = "off";
defparam \MonDReg[9]~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \MonDReg[9]~3 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_action_ocimem_a1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_b),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~2 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~2 .extended_lut = "off";
defparam \MonDReg[0]~2 .lut_mask = 64'h2727272727272727;
defparam \MonDReg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!jdo_34),
	.datad(!jdo_17),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hFF7DFFFFFF7DFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~0 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~0 .extended_lut = "off";
defparam \MonDReg~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \MonDReg~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~1 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_3),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!\MonDReg~0_combout ),
	.datae(!q_a_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~1 .extended_lut = "off";
defparam \MonDReg~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!jdo_5),
	.datae(!q_a_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_3),
	.datae(!jdo_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~6 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_4),
	.datae(!jdo_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~6 .extended_lut = "off";
defparam \MonDReg~6 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[27]~16 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[27]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[27]~16 .extended_lut = "off";
defparam \MonDReg[27]~16 .lut_mask = 64'h6666666666666666;
defparam \MonDReg[27]~16 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[27]~7 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_30),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!\MonAReg[3]~q ),
	.datae(!q_a_27),
	.dataf(!\MonDReg[27]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[27]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[27]~7 .extended_lut = "off";
defparam \MonDReg[27]~7 .lut_mask = 64'hFF7BFFFFFFFFFFFF;
defparam \MonDReg[27]~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[27]~8 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[27]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[27]~8 .extended_lut = "off";
defparam \MonDReg[27]~8 .lut_mask = 64'h2727272727272727;
defparam \MonDReg[27]~8 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~9 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_11),
	.datae(!jdo_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~9 .extended_lut = "off";
defparam \MonDReg~9 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~9 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~10 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_12),
	.datae(!jdo_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~10 .extended_lut = "off";
defparam \MonDReg~10 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~10 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~17 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~17 .extended_lut = "off";
defparam \MonDReg~17 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg~17 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~11 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_8),
	.datac(!\MonAReg[2]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_5),
	.dataf(!\MonDReg~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~11 .extended_lut = "off";
defparam \MonDReg~11 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \MonDReg~11 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[8]~12 (
	.dataa(!take_action_ocimem_b),
	.datab(!\MonAReg[2]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_8),
	.dataf(!jdo_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[8]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[8]~12 .extended_lut = "off";
defparam \MonDReg[8]~12 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \MonDReg[8]~12 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~13 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_10),
	.datae(!jdo_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~13 .extended_lut = "off";
defparam \MonDReg~13 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~13 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~19 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~19 .extended_lut = "off";
defparam \MonDReg~19 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \MonDReg~19 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~14 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_32),
	.datac(!\MonAReg[2]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_29),
	.dataf(!\MonDReg~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~14 .extended_lut = "off";
defparam \MonDReg~14 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \MonDReg~14 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~18 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~18 .extended_lut = "off";
defparam \MonDReg~18 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \MonDReg~18 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~15 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_21),
	.datac(!\MonAReg[2]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_18),
	.dataf(!\MonDReg~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~15 .extended_lut = "off";
defparam \MonDReg~15 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \MonDReg~15 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_4,
	q_a_3,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_5,
	q_a_8,
	q_a_10,
	q_a_9,
	q_a_28,
	q_a_21,
	q_a_29,
	q_a_30,
	q_a_31,
	q_a_17,
	q_a_18,
	q_a_27,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_22,
	ociram_byteenable_2,
	ociram_wr_data_23,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_4,
	ociram_wr_data_3,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_12,
	ociram_wr_data_13,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_16,
	ociram_wr_data_5,
	ociram_wr_data_8,
	ociram_wr_data_10,
	ociram_wr_data_9,
	ociram_wr_data_28,
	ociram_wr_data_21,
	ociram_wr_data_29,
	ociram_wr_data_30,
	ociram_wr_data_31,
	ociram_wr_data_17,
	ociram_wr_data_18,
	ociram_wr_data_27,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_20,
	ociram_wr_data_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_4;
output 	q_a_3;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_5;
output 	q_a_8;
output 	q_a_10;
output 	q_a_9;
output 	q_a_28;
output 	q_a_21;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	q_a_17;
output 	q_a_18;
output 	q_a_27;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_19;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_22;
input 	ociram_byteenable_2;
input 	ociram_wr_data_23;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_4;
input 	ociram_wr_data_3;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_12;
input 	ociram_wr_data_13;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_16;
input 	ociram_wr_data_5;
input 	ociram_wr_data_8;
input 	ociram_wr_data_10;
input 	ociram_wr_data_9;
input 	ociram_wr_data_28;
input 	ociram_wr_data_21;
input 	ociram_wr_data_29;
input 	ociram_wr_data_30;
input 	ociram_wr_data_31;
input 	ociram_wr_data_17;
input 	ociram_wr_data_18;
input 	ociram_wr_data_27;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module sdram_demo_altsyncram_1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[13:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_qid1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module sdram_demo_altsyncram_qid1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_nios2_oci:the_sdram_demo_nios2_cpu_nios2_oci|sdram_demo_nios2_cpu_nios2_ocimem:the_sdram_demo_nios2_cpu_nios2_ocimem|sdram_demo_nios2_cpu_ociram_sp_ram_module:sdram_demo_nios2_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_register_bank_a_module (
	q_b_4,
	q_b_5,
	q_b_9,
	D_iw_28,
	q_b_24,
	D_iw_29,
	q_b_25,
	D_iw_30,
	q_b_26,
	D_iw_31,
	q_b_27,
	q_b_28,
	q_b_20,
	q_b_19,
	q_b_21,
	q_b_22,
	D_iw_27,
	q_b_23,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_2,
	q_b_3,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_1,
	q_b_0,
	W_rf_wr_data_0,
	W_rf_wren,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_9,
	W_rf_wr_data_24,
	W_rf_wr_data_25,
	W_rf_wr_data_26,
	W_rf_wr_data_27,
	W_rf_wr_data_28,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_21,
	W_rf_wr_data_22,
	W_rf_wr_data_23,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_8,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_5;
output 	q_b_9;
input 	D_iw_28;
output 	q_b_24;
input 	D_iw_29;
output 	q_b_25;
input 	D_iw_30;
output 	q_b_26;
input 	D_iw_31;
output 	q_b_27;
output 	q_b_28;
output 	q_b_20;
output 	q_b_19;
output 	q_b_21;
output 	q_b_22;
input 	D_iw_27;
output 	q_b_23;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_2;
output 	q_b_3;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_1;
output 	q_b_0;
input 	W_rf_wr_data_0;
input 	W_rf_wren;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.wren_a(W_rf_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module sdram_demo_altsyncram_2 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[13:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_msi1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module sdram_demo_altsyncram_msi1 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_a_module:sdram_demo_nios2_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module sdram_demo_sdram_demo_nios2_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	D_iw_22,
	D_iw_23,
	D_iw_24,
	D_iw_25,
	D_iw_26,
	q_b_9,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_20,
	q_b_19,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_8,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_31,
	q_b_30,
	q_b_29,
	W_rf_wr_data_0,
	W_rf_wren,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_9,
	W_rf_wr_data_24,
	W_rf_wr_data_25,
	W_rf_wr_data_26,
	W_rf_wr_data_27,
	W_rf_wr_data_28,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_21,
	W_rf_wr_data_22,
	W_rf_wr_data_23,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_8,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	D_iw_22;
input 	D_iw_23;
input 	D_iw_24;
input 	D_iw_25;
input 	D_iw_26;
output 	q_b_9;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_20;
output 	q_b_19;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_8;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
input 	W_rf_wr_data_0;
input 	W_rf_wren;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.wren_a(W_rf_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module sdram_demo_altsyncram_3 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[13:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_msi1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module sdram_demo_altsyncram_msi1_1 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "sdram_demo_nios2:nios2|sdram_demo_nios2_cpu:cpu|sdram_demo_nios2_cpu_register_bank_b_module:sdram_demo_nios2_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module sdram_demo_sdram_demo_ram (
	ram_block1a32,
	ram_block1a0,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a37,
	ram_block1a5,
	ram_block1a40,
	ram_block1a8,
	ram_block1a42,
	ram_block1a10,
	ram_block1a41,
	ram_block1a9,
	ram_block1a60,
	ram_block1a28,
	ram_block1a53,
	ram_block1a21,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	ram_block1a52,
	ram_block1a20,
	ram_block1a51,
	ram_block1a19,
	d_write,
	write_accepted,
	saved_grant_0,
	mem_used_1,
	Equal1,
	src5_valid,
	src_valid,
	address_reg_a_0,
	r_early_rst,
	src_data_51,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_33,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a32;
output 	ram_block1a0;
output 	ram_block1a54;
output 	ram_block1a22;
output 	ram_block1a55;
output 	ram_block1a23;
output 	ram_block1a56;
output 	ram_block1a24;
output 	ram_block1a57;
output 	ram_block1a25;
output 	ram_block1a58;
output 	ram_block1a26;
output 	ram_block1a33;
output 	ram_block1a1;
output 	ram_block1a36;
output 	ram_block1a4;
output 	ram_block1a35;
output 	ram_block1a3;
output 	ram_block1a34;
output 	ram_block1a2;
output 	ram_block1a43;
output 	ram_block1a11;
output 	ram_block1a44;
output 	ram_block1a12;
output 	ram_block1a45;
output 	ram_block1a13;
output 	ram_block1a46;
output 	ram_block1a14;
output 	ram_block1a47;
output 	ram_block1a15;
output 	ram_block1a48;
output 	ram_block1a16;
output 	ram_block1a37;
output 	ram_block1a5;
output 	ram_block1a40;
output 	ram_block1a8;
output 	ram_block1a42;
output 	ram_block1a10;
output 	ram_block1a41;
output 	ram_block1a9;
output 	ram_block1a60;
output 	ram_block1a28;
output 	ram_block1a53;
output 	ram_block1a21;
output 	ram_block1a61;
output 	ram_block1a29;
output 	ram_block1a62;
output 	ram_block1a30;
output 	ram_block1a63;
output 	ram_block1a31;
output 	ram_block1a49;
output 	ram_block1a17;
output 	ram_block1a50;
output 	ram_block1a18;
output 	ram_block1a59;
output 	ram_block1a27;
output 	ram_block1a39;
output 	ram_block1a7;
output 	ram_block1a38;
output 	ram_block1a6;
output 	ram_block1a52;
output 	ram_block1a20;
output 	ram_block1a51;
output 	ram_block1a19;
input 	d_write;
input 	write_accepted;
input 	saved_grant_0;
input 	mem_used_1;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
output 	address_reg_a_0;
input 	r_early_rst;
input 	src_data_51;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_data_33;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;
wire \wren~1_combout ;


sdram_demo_altsyncram_4 the_altsyncram(
	.ram_block1a32(ram_block1a32),
	.ram_block1a0(ram_block1a0),
	.ram_block1a54(ram_block1a54),
	.ram_block1a22(ram_block1a22),
	.ram_block1a55(ram_block1a55),
	.ram_block1a23(ram_block1a23),
	.ram_block1a56(ram_block1a56),
	.ram_block1a24(ram_block1a24),
	.ram_block1a57(ram_block1a57),
	.ram_block1a25(ram_block1a25),
	.ram_block1a58(ram_block1a58),
	.ram_block1a26(ram_block1a26),
	.ram_block1a33(ram_block1a33),
	.ram_block1a1(ram_block1a1),
	.ram_block1a36(ram_block1a36),
	.ram_block1a4(ram_block1a4),
	.ram_block1a35(ram_block1a35),
	.ram_block1a3(ram_block1a3),
	.ram_block1a34(ram_block1a34),
	.ram_block1a2(ram_block1a2),
	.ram_block1a43(ram_block1a43),
	.ram_block1a11(ram_block1a11),
	.ram_block1a44(ram_block1a44),
	.ram_block1a12(ram_block1a12),
	.ram_block1a45(ram_block1a45),
	.ram_block1a13(ram_block1a13),
	.ram_block1a46(ram_block1a46),
	.ram_block1a14(ram_block1a14),
	.ram_block1a47(ram_block1a47),
	.ram_block1a15(ram_block1a15),
	.ram_block1a48(ram_block1a48),
	.ram_block1a16(ram_block1a16),
	.ram_block1a37(ram_block1a37),
	.ram_block1a5(ram_block1a5),
	.ram_block1a40(ram_block1a40),
	.ram_block1a8(ram_block1a8),
	.ram_block1a42(ram_block1a42),
	.ram_block1a10(ram_block1a10),
	.ram_block1a41(ram_block1a41),
	.ram_block1a9(ram_block1a9),
	.ram_block1a60(ram_block1a60),
	.ram_block1a28(ram_block1a28),
	.ram_block1a53(ram_block1a53),
	.ram_block1a21(ram_block1a21),
	.ram_block1a61(ram_block1a61),
	.ram_block1a29(ram_block1a29),
	.ram_block1a62(ram_block1a62),
	.ram_block1a30(ram_block1a30),
	.ram_block1a63(ram_block1a63),
	.ram_block1a31(ram_block1a31),
	.ram_block1a49(ram_block1a49),
	.ram_block1a17(ram_block1a17),
	.ram_block1a50(ram_block1a50),
	.ram_block1a18(ram_block1a18),
	.ram_block1a59(ram_block1a59),
	.ram_block1a27(ram_block1a27),
	.ram_block1a39(ram_block1a39),
	.ram_block1a7(ram_block1a7),
	.ram_block1a38(ram_block1a38),
	.ram_block1a6(ram_block1a6),
	.ram_block1a52(ram_block1a52),
	.ram_block1a20(ram_block1a20),
	.ram_block1a51(ram_block1a51),
	.ram_block1a19(ram_block1a19),
	.saved_grant_0(saved_grant_0),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.address_reg_a_0(address_reg_a_0),
	.clocken0(r_early_rst),
	.address_a({src_data_51,src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.wren(\wren~0_combout ),
	.wren1(\wren~1_combout ),
	.data_a({src_payload24,src_payload23,src_payload22,src_payload20,src_payload27,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload21,src_payload30,src_payload31,src_payload26,src_payload25,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,
src_payload10,src_payload18,src_payload19,src_payload17,src_payload28,src_payload29,src_payload16,src_payload7,src_payload8,src_payload9,src_payload6,src_payload}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!write_accepted),
	.datac(!saved_grant_0),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \wren~0 .shared_arith = "off";

cyclonev_lcell_comb \wren~1 (
	.dataa(!saved_grant_0),
	.datab(!Equal1),
	.datac(!src5_valid),
	.datad(!src_valid),
	.datae(!\wren~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~1 .extended_lut = "off";
defparam \wren~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \wren~1 .shared_arith = "off";

endmodule

module sdram_demo_altsyncram_4 (
	ram_block1a32,
	ram_block1a0,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a33,
	ram_block1a1,
	ram_block1a36,
	ram_block1a4,
	ram_block1a35,
	ram_block1a3,
	ram_block1a34,
	ram_block1a2,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a37,
	ram_block1a5,
	ram_block1a40,
	ram_block1a8,
	ram_block1a42,
	ram_block1a10,
	ram_block1a41,
	ram_block1a9,
	ram_block1a60,
	ram_block1a28,
	ram_block1a53,
	ram_block1a21,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a59,
	ram_block1a27,
	ram_block1a39,
	ram_block1a7,
	ram_block1a38,
	ram_block1a6,
	ram_block1a52,
	ram_block1a20,
	ram_block1a51,
	ram_block1a19,
	saved_grant_0,
	Equal1,
	src5_valid,
	src_valid,
	address_reg_a_0,
	clocken0,
	address_a,
	wren,
	wren1,
	data_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a32;
output 	ram_block1a0;
output 	ram_block1a54;
output 	ram_block1a22;
output 	ram_block1a55;
output 	ram_block1a23;
output 	ram_block1a56;
output 	ram_block1a24;
output 	ram_block1a57;
output 	ram_block1a25;
output 	ram_block1a58;
output 	ram_block1a26;
output 	ram_block1a33;
output 	ram_block1a1;
output 	ram_block1a36;
output 	ram_block1a4;
output 	ram_block1a35;
output 	ram_block1a3;
output 	ram_block1a34;
output 	ram_block1a2;
output 	ram_block1a43;
output 	ram_block1a11;
output 	ram_block1a44;
output 	ram_block1a12;
output 	ram_block1a45;
output 	ram_block1a13;
output 	ram_block1a46;
output 	ram_block1a14;
output 	ram_block1a47;
output 	ram_block1a15;
output 	ram_block1a48;
output 	ram_block1a16;
output 	ram_block1a37;
output 	ram_block1a5;
output 	ram_block1a40;
output 	ram_block1a8;
output 	ram_block1a42;
output 	ram_block1a10;
output 	ram_block1a41;
output 	ram_block1a9;
output 	ram_block1a60;
output 	ram_block1a28;
output 	ram_block1a53;
output 	ram_block1a21;
output 	ram_block1a61;
output 	ram_block1a29;
output 	ram_block1a62;
output 	ram_block1a30;
output 	ram_block1a63;
output 	ram_block1a31;
output 	ram_block1a49;
output 	ram_block1a17;
output 	ram_block1a50;
output 	ram_block1a18;
output 	ram_block1a59;
output 	ram_block1a27;
output 	ram_block1a39;
output 	ram_block1a7;
output 	ram_block1a38;
output 	ram_block1a6;
output 	ram_block1a52;
output 	ram_block1a20;
output 	ram_block1a51;
output 	ram_block1a19;
input 	saved_grant_0;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
output 	address_reg_a_0;
input 	clocken0;
input 	[13:0] address_a;
input 	wren;
input 	wren1;
input 	[31:0] data_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sdram_demo_altsyncram_pgm1 auto_generated(
	.ram_block1a321(ram_block1a32),
	.ram_block1a01(ram_block1a0),
	.ram_block1a541(ram_block1a54),
	.ram_block1a221(ram_block1a22),
	.ram_block1a551(ram_block1a55),
	.ram_block1a231(ram_block1a23),
	.ram_block1a561(ram_block1a56),
	.ram_block1a241(ram_block1a24),
	.ram_block1a571(ram_block1a57),
	.ram_block1a251(ram_block1a25),
	.ram_block1a581(ram_block1a58),
	.ram_block1a261(ram_block1a26),
	.ram_block1a331(ram_block1a33),
	.ram_block1a110(ram_block1a1),
	.ram_block1a361(ram_block1a36),
	.ram_block1a410(ram_block1a4),
	.ram_block1a351(ram_block1a35),
	.ram_block1a310(ram_block1a3),
	.ram_block1a341(ram_block1a34),
	.ram_block1a210(ram_block1a2),
	.ram_block1a431(ram_block1a43),
	.ram_block1a111(ram_block1a11),
	.ram_block1a441(ram_block1a44),
	.ram_block1a121(ram_block1a12),
	.ram_block1a451(ram_block1a45),
	.ram_block1a131(ram_block1a13),
	.ram_block1a461(ram_block1a46),
	.ram_block1a141(ram_block1a14),
	.ram_block1a471(ram_block1a47),
	.ram_block1a151(ram_block1a15),
	.ram_block1a481(ram_block1a48),
	.ram_block1a161(ram_block1a16),
	.ram_block1a371(ram_block1a37),
	.ram_block1a510(ram_block1a5),
	.ram_block1a401(ram_block1a40),
	.ram_block1a81(ram_block1a8),
	.ram_block1a421(ram_block1a42),
	.ram_block1a101(ram_block1a10),
	.ram_block1a411(ram_block1a41),
	.ram_block1a91(ram_block1a9),
	.ram_block1a601(ram_block1a60),
	.ram_block1a281(ram_block1a28),
	.ram_block1a531(ram_block1a53),
	.ram_block1a211(ram_block1a21),
	.ram_block1a611(ram_block1a61),
	.ram_block1a291(ram_block1a29),
	.ram_block1a621(ram_block1a62),
	.ram_block1a301(ram_block1a30),
	.ram_block1a631(ram_block1a63),
	.ram_block1a311(ram_block1a31),
	.ram_block1a491(ram_block1a49),
	.ram_block1a171(ram_block1a17),
	.ram_block1a501(ram_block1a50),
	.ram_block1a181(ram_block1a18),
	.ram_block1a591(ram_block1a59),
	.ram_block1a271(ram_block1a27),
	.ram_block1a391(ram_block1a39),
	.ram_block1a71(ram_block1a7),
	.ram_block1a381(ram_block1a38),
	.ram_block1a64(ram_block1a6),
	.ram_block1a521(ram_block1a52),
	.ram_block1a201(ram_block1a20),
	.ram_block1a511(ram_block1a51),
	.ram_block1a191(ram_block1a19),
	.saved_grant_0(saved_grant_0),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.address_reg_a_0(address_reg_a_0),
	.clocken0(clocken0),
	.address_a({address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren(wren),
	.wren1(wren1),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module sdram_demo_altsyncram_pgm1 (
	ram_block1a321,
	ram_block1a01,
	ram_block1a541,
	ram_block1a221,
	ram_block1a551,
	ram_block1a231,
	ram_block1a561,
	ram_block1a241,
	ram_block1a571,
	ram_block1a251,
	ram_block1a581,
	ram_block1a261,
	ram_block1a331,
	ram_block1a110,
	ram_block1a361,
	ram_block1a410,
	ram_block1a351,
	ram_block1a310,
	ram_block1a341,
	ram_block1a210,
	ram_block1a431,
	ram_block1a111,
	ram_block1a441,
	ram_block1a121,
	ram_block1a451,
	ram_block1a131,
	ram_block1a461,
	ram_block1a141,
	ram_block1a471,
	ram_block1a151,
	ram_block1a481,
	ram_block1a161,
	ram_block1a371,
	ram_block1a510,
	ram_block1a401,
	ram_block1a81,
	ram_block1a421,
	ram_block1a101,
	ram_block1a411,
	ram_block1a91,
	ram_block1a601,
	ram_block1a281,
	ram_block1a531,
	ram_block1a211,
	ram_block1a611,
	ram_block1a291,
	ram_block1a621,
	ram_block1a301,
	ram_block1a631,
	ram_block1a311,
	ram_block1a491,
	ram_block1a171,
	ram_block1a501,
	ram_block1a181,
	ram_block1a591,
	ram_block1a271,
	ram_block1a391,
	ram_block1a71,
	ram_block1a381,
	ram_block1a64,
	ram_block1a521,
	ram_block1a201,
	ram_block1a511,
	ram_block1a191,
	saved_grant_0,
	Equal1,
	src5_valid,
	src_valid,
	address_reg_a_0,
	clocken0,
	address_a,
	wren,
	wren1,
	data_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a321;
output 	ram_block1a01;
output 	ram_block1a541;
output 	ram_block1a221;
output 	ram_block1a551;
output 	ram_block1a231;
output 	ram_block1a561;
output 	ram_block1a241;
output 	ram_block1a571;
output 	ram_block1a251;
output 	ram_block1a581;
output 	ram_block1a261;
output 	ram_block1a331;
output 	ram_block1a110;
output 	ram_block1a361;
output 	ram_block1a410;
output 	ram_block1a351;
output 	ram_block1a310;
output 	ram_block1a341;
output 	ram_block1a210;
output 	ram_block1a431;
output 	ram_block1a111;
output 	ram_block1a441;
output 	ram_block1a121;
output 	ram_block1a451;
output 	ram_block1a131;
output 	ram_block1a461;
output 	ram_block1a141;
output 	ram_block1a471;
output 	ram_block1a151;
output 	ram_block1a481;
output 	ram_block1a161;
output 	ram_block1a371;
output 	ram_block1a510;
output 	ram_block1a401;
output 	ram_block1a81;
output 	ram_block1a421;
output 	ram_block1a101;
output 	ram_block1a411;
output 	ram_block1a91;
output 	ram_block1a601;
output 	ram_block1a281;
output 	ram_block1a531;
output 	ram_block1a211;
output 	ram_block1a611;
output 	ram_block1a291;
output 	ram_block1a621;
output 	ram_block1a301;
output 	ram_block1a631;
output 	ram_block1a311;
output 	ram_block1a491;
output 	ram_block1a171;
output 	ram_block1a501;
output 	ram_block1a181;
output 	ram_block1a591;
output 	ram_block1a271;
output 	ram_block1a391;
output 	ram_block1a71;
output 	ram_block1a381;
output 	ram_block1a64;
output 	ram_block1a521;
output 	ram_block1a201;
output 	ram_block1a511;
output 	ram_block1a191;
input 	saved_grant_0;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
output 	address_reg_a_0;
input 	clocken0;
input 	[13:0] address_a;
input 	wren;
input 	wren1;
input 	[31:0] data_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \decode3|eq_node[1]~combout ;
wire \decode3|eq_node[0]~combout ;

wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;

assign ram_block1a321 = ram_block1a32_PORTADATAOUT_bus[0];

assign ram_block1a01 = ram_block1a0_PORTADATAOUT_bus[0];

assign ram_block1a541 = ram_block1a54_PORTADATAOUT_bus[0];

assign ram_block1a221 = ram_block1a22_PORTADATAOUT_bus[0];

assign ram_block1a551 = ram_block1a55_PORTADATAOUT_bus[0];

assign ram_block1a231 = ram_block1a23_PORTADATAOUT_bus[0];

assign ram_block1a561 = ram_block1a56_PORTADATAOUT_bus[0];

assign ram_block1a241 = ram_block1a24_PORTADATAOUT_bus[0];

assign ram_block1a571 = ram_block1a57_PORTADATAOUT_bus[0];

assign ram_block1a251 = ram_block1a25_PORTADATAOUT_bus[0];

assign ram_block1a581 = ram_block1a58_PORTADATAOUT_bus[0];

assign ram_block1a261 = ram_block1a26_PORTADATAOUT_bus[0];

assign ram_block1a331 = ram_block1a33_PORTADATAOUT_bus[0];

assign ram_block1a110 = ram_block1a1_PORTADATAOUT_bus[0];

assign ram_block1a361 = ram_block1a36_PORTADATAOUT_bus[0];

assign ram_block1a410 = ram_block1a4_PORTADATAOUT_bus[0];

assign ram_block1a351 = ram_block1a35_PORTADATAOUT_bus[0];

assign ram_block1a310 = ram_block1a3_PORTADATAOUT_bus[0];

assign ram_block1a341 = ram_block1a34_PORTADATAOUT_bus[0];

assign ram_block1a210 = ram_block1a2_PORTADATAOUT_bus[0];

assign ram_block1a431 = ram_block1a43_PORTADATAOUT_bus[0];

assign ram_block1a111 = ram_block1a11_PORTADATAOUT_bus[0];

assign ram_block1a441 = ram_block1a44_PORTADATAOUT_bus[0];

assign ram_block1a121 = ram_block1a12_PORTADATAOUT_bus[0];

assign ram_block1a451 = ram_block1a45_PORTADATAOUT_bus[0];

assign ram_block1a131 = ram_block1a13_PORTADATAOUT_bus[0];

assign ram_block1a461 = ram_block1a46_PORTADATAOUT_bus[0];

assign ram_block1a141 = ram_block1a14_PORTADATAOUT_bus[0];

assign ram_block1a471 = ram_block1a47_PORTADATAOUT_bus[0];

assign ram_block1a151 = ram_block1a15_PORTADATAOUT_bus[0];

assign ram_block1a481 = ram_block1a48_PORTADATAOUT_bus[0];

assign ram_block1a161 = ram_block1a16_PORTADATAOUT_bus[0];

assign ram_block1a371 = ram_block1a37_PORTADATAOUT_bus[0];

assign ram_block1a510 = ram_block1a5_PORTADATAOUT_bus[0];

assign ram_block1a401 = ram_block1a40_PORTADATAOUT_bus[0];

assign ram_block1a81 = ram_block1a8_PORTADATAOUT_bus[0];

assign ram_block1a421 = ram_block1a42_PORTADATAOUT_bus[0];

assign ram_block1a101 = ram_block1a10_PORTADATAOUT_bus[0];

assign ram_block1a411 = ram_block1a41_PORTADATAOUT_bus[0];

assign ram_block1a91 = ram_block1a9_PORTADATAOUT_bus[0];

assign ram_block1a601 = ram_block1a60_PORTADATAOUT_bus[0];

assign ram_block1a281 = ram_block1a28_PORTADATAOUT_bus[0];

assign ram_block1a531 = ram_block1a53_PORTADATAOUT_bus[0];

assign ram_block1a211 = ram_block1a21_PORTADATAOUT_bus[0];

assign ram_block1a611 = ram_block1a61_PORTADATAOUT_bus[0];

assign ram_block1a291 = ram_block1a29_PORTADATAOUT_bus[0];

assign ram_block1a621 = ram_block1a62_PORTADATAOUT_bus[0];

assign ram_block1a301 = ram_block1a30_PORTADATAOUT_bus[0];

assign ram_block1a631 = ram_block1a63_PORTADATAOUT_bus[0];

assign ram_block1a311 = ram_block1a31_PORTADATAOUT_bus[0];

assign ram_block1a491 = ram_block1a49_PORTADATAOUT_bus[0];

assign ram_block1a171 = ram_block1a17_PORTADATAOUT_bus[0];

assign ram_block1a501 = ram_block1a50_PORTADATAOUT_bus[0];

assign ram_block1a181 = ram_block1a18_PORTADATAOUT_bus[0];

assign ram_block1a591 = ram_block1a59_PORTADATAOUT_bus[0];

assign ram_block1a271 = ram_block1a27_PORTADATAOUT_bus[0];

assign ram_block1a391 = ram_block1a39_PORTADATAOUT_bus[0];

assign ram_block1a71 = ram_block1a7_PORTADATAOUT_bus[0];

assign ram_block1a381 = ram_block1a38_PORTADATAOUT_bus[0];

assign ram_block1a64 = ram_block1a6_PORTADATAOUT_bus[0];

assign ram_block1a521 = ram_block1a52_PORTADATAOUT_bus[0];

assign ram_block1a201 = ram_block1a20_PORTADATAOUT_bus[0];

assign ram_block1a511 = ram_block1a51_PORTADATAOUT_bus[0];

assign ram_block1a191 = ram_block1a19_PORTADATAOUT_bus[0];

sdram_demo_decode_5la decode3(
	.saved_grant_0(saved_grant_0),
	.Equal1(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.src_data_51(address_a[13]),
	.wren(wren),
	.eq_node_1(\decode3|eq_node[1]~combout ),
	.eq_node_0(\decode3|eq_node[0]~combout ));

cyclonev_ram_block ram_block1a32(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.init_file = "sdram_demo_ram.hex";
defparam ram_block1a32.init_file_layout = "port_a";
defparam ram_block1a32.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.operation_mode = "single_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_byte_enable_mask_width = 1;
defparam ram_block1a32.port_a_byte_size = 1;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 8192;
defparam ram_block1a32.port_a_first_bit_number = 0;
defparam ram_block1a32.port_a_last_address = 16383;
defparam ram_block1a32.port_a_logical_ram_depth = 16384;
defparam ram_block1a32.port_a_logical_ram_width = 32;
defparam ram_block1a32.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a32.ram_block_type = "auto";
defparam ram_block1a32.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a32.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a32.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a32.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a0(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "sdram_demo_ram.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 16384;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a54(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.init_file = "sdram_demo_ram.hex";
defparam ram_block1a54.init_file_layout = "port_a";
defparam ram_block1a54.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.operation_mode = "single_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_byte_enable_mask_width = 1;
defparam ram_block1a54.port_a_byte_size = 1;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 8192;
defparam ram_block1a54.port_a_first_bit_number = 22;
defparam ram_block1a54.port_a_last_address = 16383;
defparam ram_block1a54.port_a_logical_ram_depth = 16384;
defparam ram_block1a54.port_a_logical_ram_width = 32;
defparam ram_block1a54.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a54.ram_block_type = "auto";
defparam ram_block1a54.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a54.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a54.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a54.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "sdram_demo_ram.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 16384;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a55(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.init_file = "sdram_demo_ram.hex";
defparam ram_block1a55.init_file_layout = "port_a";
defparam ram_block1a55.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.operation_mode = "single_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_byte_enable_mask_width = 1;
defparam ram_block1a55.port_a_byte_size = 1;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 8192;
defparam ram_block1a55.port_a_first_bit_number = 23;
defparam ram_block1a55.port_a_last_address = 16383;
defparam ram_block1a55.port_a_logical_ram_depth = 16384;
defparam ram_block1a55.port_a_logical_ram_width = 32;
defparam ram_block1a55.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a55.ram_block_type = "auto";
defparam ram_block1a55.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a55.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a55.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a55.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "sdram_demo_ram.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 16384;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a56(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.init_file = "sdram_demo_ram.hex";
defparam ram_block1a56.init_file_layout = "port_a";
defparam ram_block1a56.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.operation_mode = "single_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_byte_enable_mask_width = 1;
defparam ram_block1a56.port_a_byte_size = 1;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 8192;
defparam ram_block1a56.port_a_first_bit_number = 24;
defparam ram_block1a56.port_a_last_address = 16383;
defparam ram_block1a56.port_a_logical_ram_depth = 16384;
defparam ram_block1a56.port_a_logical_ram_width = 32;
defparam ram_block1a56.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a56.ram_block_type = "auto";
defparam ram_block1a56.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a56.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a56.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a56.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "sdram_demo_ram.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 16384;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a57(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.init_file = "sdram_demo_ram.hex";
defparam ram_block1a57.init_file_layout = "port_a";
defparam ram_block1a57.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.operation_mode = "single_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_byte_enable_mask_width = 1;
defparam ram_block1a57.port_a_byte_size = 1;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 8192;
defparam ram_block1a57.port_a_first_bit_number = 25;
defparam ram_block1a57.port_a_last_address = 16383;
defparam ram_block1a57.port_a_logical_ram_depth = 16384;
defparam ram_block1a57.port_a_logical_ram_width = 32;
defparam ram_block1a57.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a57.ram_block_type = "auto";
defparam ram_block1a57.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a57.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a57.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a57.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "sdram_demo_ram.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 16384;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a58(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.init_file = "sdram_demo_ram.hex";
defparam ram_block1a58.init_file_layout = "port_a";
defparam ram_block1a58.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.operation_mode = "single_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_byte_enable_mask_width = 1;
defparam ram_block1a58.port_a_byte_size = 1;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 8192;
defparam ram_block1a58.port_a_first_bit_number = 26;
defparam ram_block1a58.port_a_last_address = 16383;
defparam ram_block1a58.port_a_logical_ram_depth = 16384;
defparam ram_block1a58.port_a_logical_ram_width = 32;
defparam ram_block1a58.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a58.ram_block_type = "auto";
defparam ram_block1a58.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a58.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a58.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a58.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "sdram_demo_ram.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 16384;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a33(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.init_file = "sdram_demo_ram.hex";
defparam ram_block1a33.init_file_layout = "port_a";
defparam ram_block1a33.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.operation_mode = "single_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_byte_enable_mask_width = 1;
defparam ram_block1a33.port_a_byte_size = 1;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 8192;
defparam ram_block1a33.port_a_first_bit_number = 1;
defparam ram_block1a33.port_a_last_address = 16383;
defparam ram_block1a33.port_a_logical_ram_depth = 16384;
defparam ram_block1a33.port_a_logical_ram_width = 32;
defparam ram_block1a33.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a33.ram_block_type = "auto";
defparam ram_block1a33.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a33.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a33.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a33.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "sdram_demo_ram.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 16384;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a36(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.init_file = "sdram_demo_ram.hex";
defparam ram_block1a36.init_file_layout = "port_a";
defparam ram_block1a36.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.operation_mode = "single_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_byte_enable_mask_width = 1;
defparam ram_block1a36.port_a_byte_size = 1;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 8192;
defparam ram_block1a36.port_a_first_bit_number = 4;
defparam ram_block1a36.port_a_last_address = 16383;
defparam ram_block1a36.port_a_logical_ram_depth = 16384;
defparam ram_block1a36.port_a_logical_ram_width = 32;
defparam ram_block1a36.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a36.ram_block_type = "auto";
defparam ram_block1a36.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a36.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a36.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a36.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a4(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "sdram_demo_ram.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 16384;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a35(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.init_file = "sdram_demo_ram.hex";
defparam ram_block1a35.init_file_layout = "port_a";
defparam ram_block1a35.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.operation_mode = "single_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_byte_enable_mask_width = 1;
defparam ram_block1a35.port_a_byte_size = 1;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 8192;
defparam ram_block1a35.port_a_first_bit_number = 3;
defparam ram_block1a35.port_a_last_address = 16383;
defparam ram_block1a35.port_a_logical_ram_depth = 16384;
defparam ram_block1a35.port_a_logical_ram_width = 32;
defparam ram_block1a35.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a35.ram_block_type = "auto";
defparam ram_block1a35.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a35.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a35.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a35.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "sdram_demo_ram.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 16384;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a34(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.init_file = "sdram_demo_ram.hex";
defparam ram_block1a34.init_file_layout = "port_a";
defparam ram_block1a34.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.operation_mode = "single_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_byte_enable_mask_width = 1;
defparam ram_block1a34.port_a_byte_size = 1;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 8192;
defparam ram_block1a34.port_a_first_bit_number = 2;
defparam ram_block1a34.port_a_last_address = 16383;
defparam ram_block1a34.port_a_logical_ram_depth = 16384;
defparam ram_block1a34.port_a_logical_ram_width = 32;
defparam ram_block1a34.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a34.ram_block_type = "auto";
defparam ram_block1a34.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a34.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a34.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a34.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "sdram_demo_ram.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 16384;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a43(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.init_file = "sdram_demo_ram.hex";
defparam ram_block1a43.init_file_layout = "port_a";
defparam ram_block1a43.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.operation_mode = "single_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_byte_enable_mask_width = 1;
defparam ram_block1a43.port_a_byte_size = 1;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 8192;
defparam ram_block1a43.port_a_first_bit_number = 11;
defparam ram_block1a43.port_a_last_address = 16383;
defparam ram_block1a43.port_a_logical_ram_depth = 16384;
defparam ram_block1a43.port_a_logical_ram_width = 32;
defparam ram_block1a43.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a43.ram_block_type = "auto";
defparam ram_block1a43.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "sdram_demo_ram.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 16384;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a44(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.init_file = "sdram_demo_ram.hex";
defparam ram_block1a44.init_file_layout = "port_a";
defparam ram_block1a44.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.operation_mode = "single_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_byte_enable_mask_width = 1;
defparam ram_block1a44.port_a_byte_size = 1;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 8192;
defparam ram_block1a44.port_a_first_bit_number = 12;
defparam ram_block1a44.port_a_last_address = 16383;
defparam ram_block1a44.port_a_logical_ram_depth = 16384;
defparam ram_block1a44.port_a_logical_ram_width = 32;
defparam ram_block1a44.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a44.ram_block_type = "auto";
defparam ram_block1a44.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "sdram_demo_ram.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 16384;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a45(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.init_file = "sdram_demo_ram.hex";
defparam ram_block1a45.init_file_layout = "port_a";
defparam ram_block1a45.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.operation_mode = "single_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_byte_enable_mask_width = 1;
defparam ram_block1a45.port_a_byte_size = 1;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 8192;
defparam ram_block1a45.port_a_first_bit_number = 13;
defparam ram_block1a45.port_a_last_address = 16383;
defparam ram_block1a45.port_a_logical_ram_depth = 16384;
defparam ram_block1a45.port_a_logical_ram_width = 32;
defparam ram_block1a45.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a45.ram_block_type = "auto";
defparam ram_block1a45.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a45.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a45.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a45.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "sdram_demo_ram.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 16384;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a46(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.init_file = "sdram_demo_ram.hex";
defparam ram_block1a46.init_file_layout = "port_a";
defparam ram_block1a46.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.operation_mode = "single_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_byte_enable_mask_width = 1;
defparam ram_block1a46.port_a_byte_size = 1;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 8192;
defparam ram_block1a46.port_a_first_bit_number = 14;
defparam ram_block1a46.port_a_last_address = 16383;
defparam ram_block1a46.port_a_logical_ram_depth = 16384;
defparam ram_block1a46.port_a_logical_ram_width = 32;
defparam ram_block1a46.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a46.ram_block_type = "auto";
defparam ram_block1a46.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a46.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a46.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a46.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "sdram_demo_ram.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 16384;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a47(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.init_file = "sdram_demo_ram.hex";
defparam ram_block1a47.init_file_layout = "port_a";
defparam ram_block1a47.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.operation_mode = "single_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_byte_enable_mask_width = 1;
defparam ram_block1a47.port_a_byte_size = 1;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 8192;
defparam ram_block1a47.port_a_first_bit_number = 15;
defparam ram_block1a47.port_a_last_address = 16383;
defparam ram_block1a47.port_a_logical_ram_depth = 16384;
defparam ram_block1a47.port_a_logical_ram_width = 32;
defparam ram_block1a47.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a47.ram_block_type = "auto";
defparam ram_block1a47.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "sdram_demo_ram.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 16384;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a48(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.init_file = "sdram_demo_ram.hex";
defparam ram_block1a48.init_file_layout = "port_a";
defparam ram_block1a48.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.operation_mode = "single_port";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_byte_enable_mask_width = 1;
defparam ram_block1a48.port_a_byte_size = 1;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "none";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 8192;
defparam ram_block1a48.port_a_first_bit_number = 16;
defparam ram_block1a48.port_a_last_address = 16383;
defparam ram_block1a48.port_a_logical_ram_depth = 16384;
defparam ram_block1a48.port_a_logical_ram_width = 32;
defparam ram_block1a48.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a48.ram_block_type = "auto";
defparam ram_block1a48.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a48.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a48.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a48.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "sdram_demo_ram.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 16384;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a37(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.init_file = "sdram_demo_ram.hex";
defparam ram_block1a37.init_file_layout = "port_a";
defparam ram_block1a37.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.operation_mode = "single_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_byte_enable_mask_width = 1;
defparam ram_block1a37.port_a_byte_size = 1;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 8192;
defparam ram_block1a37.port_a_first_bit_number = 5;
defparam ram_block1a37.port_a_last_address = 16383;
defparam ram_block1a37.port_a_logical_ram_depth = 16384;
defparam ram_block1a37.port_a_logical_ram_width = 32;
defparam ram_block1a37.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a37.ram_block_type = "auto";
defparam ram_block1a37.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a37.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a37.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a37.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "sdram_demo_ram.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 16384;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a40(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.init_file = "sdram_demo_ram.hex";
defparam ram_block1a40.init_file_layout = "port_a";
defparam ram_block1a40.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.operation_mode = "single_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_byte_enable_mask_width = 1;
defparam ram_block1a40.port_a_byte_size = 1;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 8192;
defparam ram_block1a40.port_a_first_bit_number = 8;
defparam ram_block1a40.port_a_last_address = 16383;
defparam ram_block1a40.port_a_logical_ram_depth = 16384;
defparam ram_block1a40.port_a_logical_ram_width = 32;
defparam ram_block1a40.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a40.ram_block_type = "auto";
defparam ram_block1a40.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a40.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a40.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a40.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "sdram_demo_ram.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 16384;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a42(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.init_file = "sdram_demo_ram.hex";
defparam ram_block1a42.init_file_layout = "port_a";
defparam ram_block1a42.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.operation_mode = "single_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_byte_enable_mask_width = 1;
defparam ram_block1a42.port_a_byte_size = 1;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 8192;
defparam ram_block1a42.port_a_first_bit_number = 10;
defparam ram_block1a42.port_a_last_address = 16383;
defparam ram_block1a42.port_a_logical_ram_depth = 16384;
defparam ram_block1a42.port_a_logical_ram_width = 32;
defparam ram_block1a42.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a42.ram_block_type = "auto";
defparam ram_block1a42.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a42.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a42.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a42.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "sdram_demo_ram.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 16384;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a41(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.init_file = "sdram_demo_ram.hex";
defparam ram_block1a41.init_file_layout = "port_a";
defparam ram_block1a41.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.operation_mode = "single_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_byte_enable_mask_width = 1;
defparam ram_block1a41.port_a_byte_size = 1;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 8192;
defparam ram_block1a41.port_a_first_bit_number = 9;
defparam ram_block1a41.port_a_last_address = 16383;
defparam ram_block1a41.port_a_logical_ram_depth = 16384;
defparam ram_block1a41.port_a_logical_ram_width = 32;
defparam ram_block1a41.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a41.ram_block_type = "auto";
defparam ram_block1a41.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a41.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a41.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a41.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "sdram_demo_ram.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 16384;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a60(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.init_file = "sdram_demo_ram.hex";
defparam ram_block1a60.init_file_layout = "port_a";
defparam ram_block1a60.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.operation_mode = "single_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_byte_enable_mask_width = 1;
defparam ram_block1a60.port_a_byte_size = 1;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 8192;
defparam ram_block1a60.port_a_first_bit_number = 28;
defparam ram_block1a60.port_a_last_address = 16383;
defparam ram_block1a60.port_a_logical_ram_depth = 16384;
defparam ram_block1a60.port_a_logical_ram_width = 32;
defparam ram_block1a60.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a60.ram_block_type = "auto";
defparam ram_block1a60.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "sdram_demo_ram.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 16384;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a53(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.init_file = "sdram_demo_ram.hex";
defparam ram_block1a53.init_file_layout = "port_a";
defparam ram_block1a53.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.operation_mode = "single_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_byte_enable_mask_width = 1;
defparam ram_block1a53.port_a_byte_size = 1;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 8192;
defparam ram_block1a53.port_a_first_bit_number = 21;
defparam ram_block1a53.port_a_last_address = 16383;
defparam ram_block1a53.port_a_logical_ram_depth = 16384;
defparam ram_block1a53.port_a_logical_ram_width = 32;
defparam ram_block1a53.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a53.ram_block_type = "auto";
defparam ram_block1a53.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a53.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a53.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a53.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "sdram_demo_ram.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 16384;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a61(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.init_file = "sdram_demo_ram.hex";
defparam ram_block1a61.init_file_layout = "port_a";
defparam ram_block1a61.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.operation_mode = "single_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_byte_enable_mask_width = 1;
defparam ram_block1a61.port_a_byte_size = 1;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 8192;
defparam ram_block1a61.port_a_first_bit_number = 29;
defparam ram_block1a61.port_a_last_address = 16383;
defparam ram_block1a61.port_a_logical_ram_depth = 16384;
defparam ram_block1a61.port_a_logical_ram_width = 32;
defparam ram_block1a61.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a61.ram_block_type = "auto";
defparam ram_block1a61.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "sdram_demo_ram.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 16384;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a62(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.init_file = "sdram_demo_ram.hex";
defparam ram_block1a62.init_file_layout = "port_a";
defparam ram_block1a62.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.operation_mode = "single_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_byte_enable_mask_width = 1;
defparam ram_block1a62.port_a_byte_size = 1;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 8192;
defparam ram_block1a62.port_a_first_bit_number = 30;
defparam ram_block1a62.port_a_last_address = 16383;
defparam ram_block1a62.port_a_logical_ram_depth = 16384;
defparam ram_block1a62.port_a_logical_ram_width = 32;
defparam ram_block1a62.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a62.ram_block_type = "auto";
defparam ram_block1a62.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "sdram_demo_ram.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 16384;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a63(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.init_file = "sdram_demo_ram.hex";
defparam ram_block1a63.init_file_layout = "port_a";
defparam ram_block1a63.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.operation_mode = "single_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_byte_enable_mask_width = 1;
defparam ram_block1a63.port_a_byte_size = 1;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 8192;
defparam ram_block1a63.port_a_first_bit_number = 31;
defparam ram_block1a63.port_a_last_address = 16383;
defparam ram_block1a63.port_a_logical_ram_depth = 16384;
defparam ram_block1a63.port_a_logical_ram_width = 32;
defparam ram_block1a63.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a63.ram_block_type = "auto";
defparam ram_block1a63.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "sdram_demo_ram.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 16384;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a49(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.init_file = "sdram_demo_ram.hex";
defparam ram_block1a49.init_file_layout = "port_a";
defparam ram_block1a49.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.operation_mode = "single_port";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_byte_enable_mask_width = 1;
defparam ram_block1a49.port_a_byte_size = 1;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "none";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 8192;
defparam ram_block1a49.port_a_first_bit_number = 17;
defparam ram_block1a49.port_a_last_address = 16383;
defparam ram_block1a49.port_a_logical_ram_depth = 16384;
defparam ram_block1a49.port_a_logical_ram_width = 32;
defparam ram_block1a49.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a49.ram_block_type = "auto";
defparam ram_block1a49.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a49.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a49.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a49.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "sdram_demo_ram.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 16384;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a50(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.init_file = "sdram_demo_ram.hex";
defparam ram_block1a50.init_file_layout = "port_a";
defparam ram_block1a50.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.operation_mode = "single_port";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_byte_enable_mask_width = 1;
defparam ram_block1a50.port_a_byte_size = 1;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "none";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 8192;
defparam ram_block1a50.port_a_first_bit_number = 18;
defparam ram_block1a50.port_a_last_address = 16383;
defparam ram_block1a50.port_a_logical_ram_depth = 16384;
defparam ram_block1a50.port_a_logical_ram_width = 32;
defparam ram_block1a50.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a50.ram_block_type = "auto";
defparam ram_block1a50.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a50.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a50.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a50.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "sdram_demo_ram.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 16384;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a59(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.init_file = "sdram_demo_ram.hex";
defparam ram_block1a59.init_file_layout = "port_a";
defparam ram_block1a59.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.operation_mode = "single_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_byte_enable_mask_width = 1;
defparam ram_block1a59.port_a_byte_size = 1;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 8192;
defparam ram_block1a59.port_a_first_bit_number = 27;
defparam ram_block1a59.port_a_last_address = 16383;
defparam ram_block1a59.port_a_logical_ram_depth = 16384;
defparam ram_block1a59.port_a_logical_ram_width = 32;
defparam ram_block1a59.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a59.ram_block_type = "auto";
defparam ram_block1a59.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "sdram_demo_ram.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 16384;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a39(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.init_file = "sdram_demo_ram.hex";
defparam ram_block1a39.init_file_layout = "port_a";
defparam ram_block1a39.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.operation_mode = "single_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_byte_enable_mask_width = 1;
defparam ram_block1a39.port_a_byte_size = 1;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 8192;
defparam ram_block1a39.port_a_first_bit_number = 7;
defparam ram_block1a39.port_a_last_address = 16383;
defparam ram_block1a39.port_a_logical_ram_depth = 16384;
defparam ram_block1a39.port_a_logical_ram_width = 32;
defparam ram_block1a39.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a39.ram_block_type = "auto";
defparam ram_block1a39.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a39.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a39.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a39.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "sdram_demo_ram.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 16384;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a38(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.init_file = "sdram_demo_ram.hex";
defparam ram_block1a38.init_file_layout = "port_a";
defparam ram_block1a38.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.operation_mode = "single_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_byte_enable_mask_width = 1;
defparam ram_block1a38.port_a_byte_size = 1;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 8192;
defparam ram_block1a38.port_a_first_bit_number = 6;
defparam ram_block1a38.port_a_last_address = 16383;
defparam ram_block1a38.port_a_logical_ram_depth = 16384;
defparam ram_block1a38.port_a_logical_ram_width = 32;
defparam ram_block1a38.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a38.ram_block_type = "auto";
defparam ram_block1a38.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a38.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a38.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a38.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "sdram_demo_ram.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 16384;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a52(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.init_file = "sdram_demo_ram.hex";
defparam ram_block1a52.init_file_layout = "port_a";
defparam ram_block1a52.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.operation_mode = "single_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_byte_enable_mask_width = 1;
defparam ram_block1a52.port_a_byte_size = 1;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 8192;
defparam ram_block1a52.port_a_first_bit_number = 20;
defparam ram_block1a52.port_a_last_address = 16383;
defparam ram_block1a52.port_a_logical_ram_depth = 16384;
defparam ram_block1a52.port_a_logical_ram_width = 32;
defparam ram_block1a52.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a52.ram_block_type = "auto";
defparam ram_block1a52.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a52.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a52.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a52.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "sdram_demo_ram.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 16384;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a51(
	.portawe(\decode3|eq_node[1]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.init_file = "sdram_demo_ram.hex";
defparam ram_block1a51.init_file_layout = "port_a";
defparam ram_block1a51.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.operation_mode = "single_port";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_byte_enable_mask_width = 1;
defparam ram_block1a51.port_a_byte_size = 1;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "none";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 8192;
defparam ram_block1a51.port_a_first_bit_number = 19;
defparam ram_block1a51.port_a_last_address = 16383;
defparam ram_block1a51.port_a_logical_ram_depth = 16384;
defparam ram_block1a51.port_a_logical_ram_width = 32;
defparam ram_block1a51.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a51.ram_block_type = "auto";
defparam ram_block1a51.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a51.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a51.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a51.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(\decode3|eq_node[0]~combout ),
	.portare(wren1),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "sdram_demo_ram.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "sdram_demo_ram:ram|altsyncram:the_altsyncram|altsyncram_pgm1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 16384;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clocken0),
	.q(address_reg_a_0),
	.prn(vcc));
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";

endmodule

module sdram_demo_decode_5la (
	saved_grant_0,
	Equal1,
	src5_valid,
	src_valid,
	src_data_51,
	wren,
	eq_node_1,
	eq_node_0)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_0;
input 	Equal1;
input 	src5_valid;
input 	src_valid;
input 	src_data_51;
input 	wren;
output 	eq_node_1;
output 	eq_node_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \eq_node[1] (
	.dataa(!saved_grant_0),
	.datab(!Equal1),
	.datac(!src5_valid),
	.datad(!src_valid),
	.datae(!src_data_51),
	.dataf(!wren),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[1] .extended_lut = "off";
defparam \eq_node[1] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \eq_node[1] .shared_arith = "off";

cyclonev_lcell_comb \eq_node[0] (
	.dataa(!saved_grant_0),
	.datab(!Equal1),
	.datac(!src5_valid),
	.datad(!src_valid),
	.datae(!src_data_51),
	.dataf(!wren),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[0] .extended_lut = "off";
defparam \eq_node[0] .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \eq_node[0] .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_sdram (
	m_addr_0,
	m_addr_1,
	m_addr_2,
	m_addr_3,
	m_addr_6,
	m_addr_7,
	m_addr_8,
	m_addr_9,
	oe1,
	m_addr_4,
	m_addr_5,
	m_addr_10,
	m_addr_11,
	m_addr_12,
	m_bank_0,
	m_bank_1,
	m_cmd_1,
	m_cmd_3,
	m_dqm_0,
	m_dqm_1,
	m_dqm_2,
	m_dqm_3,
	m_cmd_2,
	m_cmd_0,
	r_sync_rst,
	always0,
	entries_1,
	entries_0,
	saved_grant_0,
	WideOr0,
	za_valid1,
	Equal1,
	src5_valid,
	saved_grant_1,
	src_valid,
	src_data_68,
	src_data_58,
	src_valid1,
	src_data_59,
	src_data_60,
	src_data_61,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_50,
	src_data_51,
	m0_write,
	m0_write1,
	src_data_52,
	src_data_53,
	src_data_54,
	src_data_55,
	src_data_56,
	src_data_57,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	m_data_0,
	m_data_1,
	m_data_2,
	m_data_3,
	m_data_4,
	m_data_5,
	m_data_6,
	m_data_7,
	m_data_8,
	m_data_9,
	m_data_10,
	m_data_11,
	m_data_12,
	m_data_13,
	m_data_14,
	m_data_15,
	m_data_16,
	m_data_17,
	m_data_18,
	m_data_19,
	m_data_20,
	m_data_21,
	m_data_22,
	m_data_23,
	m_data_24,
	m_data_25,
	m_data_26,
	m_data_27,
	m_data_28,
	m_data_29,
	m_data_30,
	m_data_31,
	za_data_0,
	za_data_22,
	za_data_23,
	za_data_24,
	za_data_25,
	za_data_26,
	za_data_1,
	za_data_4,
	za_data_3,
	za_data_2,
	za_data_11,
	za_data_12,
	za_data_13,
	za_data_14,
	za_data_15,
	za_data_16,
	za_data_5,
	za_data_8,
	za_data_10,
	za_data_9,
	za_data_28,
	za_data_21,
	za_data_29,
	za_data_30,
	za_data_31,
	za_data_17,
	za_data_18,
	za_data_27,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_19,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	sdram_wire_dq_0,
	sdram_wire_dq_1,
	sdram_wire_dq_2,
	sdram_wire_dq_3,
	sdram_wire_dq_4,
	sdram_wire_dq_5,
	sdram_wire_dq_6,
	sdram_wire_dq_7,
	sdram_wire_dq_8,
	sdram_wire_dq_9,
	sdram_wire_dq_10,
	sdram_wire_dq_11,
	sdram_wire_dq_12,
	sdram_wire_dq_13,
	sdram_wire_dq_14,
	sdram_wire_dq_15,
	sdram_wire_dq_16,
	sdram_wire_dq_17,
	sdram_wire_dq_18,
	sdram_wire_dq_19,
	sdram_wire_dq_20,
	sdram_wire_dq_21,
	sdram_wire_dq_22,
	sdram_wire_dq_23,
	sdram_wire_dq_24,
	sdram_wire_dq_25,
	sdram_wire_dq_26,
	sdram_wire_dq_27,
	sdram_wire_dq_28,
	sdram_wire_dq_29,
	sdram_wire_dq_30,
	sdram_wire_dq_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	m_addr_0;
output 	m_addr_1;
output 	m_addr_2;
output 	m_addr_3;
output 	m_addr_6;
output 	m_addr_7;
output 	m_addr_8;
output 	m_addr_9;
output 	oe1;
output 	m_addr_4;
output 	m_addr_5;
output 	m_addr_10;
output 	m_addr_11;
output 	m_addr_12;
output 	m_bank_0;
output 	m_bank_1;
output 	m_cmd_1;
output 	m_cmd_3;
output 	m_dqm_0;
output 	m_dqm_1;
output 	m_dqm_2;
output 	m_dqm_3;
output 	m_cmd_2;
output 	m_cmd_0;
input 	r_sync_rst;
input 	always0;
output 	entries_1;
output 	entries_0;
input 	saved_grant_0;
input 	WideOr0;
output 	za_valid1;
input 	Equal1;
input 	src5_valid;
input 	saved_grant_1;
input 	src_valid;
input 	src_data_68;
input 	src_data_58;
input 	src_valid1;
input 	src_data_59;
input 	src_data_60;
input 	src_data_61;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
input 	src_data_50;
input 	src_data_51;
input 	m0_write;
input 	m0_write1;
input 	src_data_52;
input 	src_data_53;
input 	src_data_54;
input 	src_data_55;
input 	src_data_56;
input 	src_data_57;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	m_data_0;
output 	m_data_1;
output 	m_data_2;
output 	m_data_3;
output 	m_data_4;
output 	m_data_5;
output 	m_data_6;
output 	m_data_7;
output 	m_data_8;
output 	m_data_9;
output 	m_data_10;
output 	m_data_11;
output 	m_data_12;
output 	m_data_13;
output 	m_data_14;
output 	m_data_15;
output 	m_data_16;
output 	m_data_17;
output 	m_data_18;
output 	m_data_19;
output 	m_data_20;
output 	m_data_21;
output 	m_data_22;
output 	m_data_23;
output 	m_data_24;
output 	m_data_25;
output 	m_data_26;
output 	m_data_27;
output 	m_data_28;
output 	m_data_29;
output 	m_data_30;
output 	m_data_31;
output 	za_data_0;
output 	za_data_22;
output 	za_data_23;
output 	za_data_24;
output 	za_data_25;
output 	za_data_26;
output 	za_data_1;
output 	za_data_4;
output 	za_data_3;
output 	za_data_2;
output 	za_data_11;
output 	za_data_12;
output 	za_data_13;
output 	za_data_14;
output 	za_data_15;
output 	za_data_16;
output 	za_data_5;
output 	za_data_8;
output 	za_data_10;
output 	za_data_9;
output 	za_data_28;
output 	za_data_21;
output 	za_data_29;
output 	za_data_30;
output 	za_data_31;
output 	za_data_17;
output 	za_data_18;
output 	za_data_27;
output 	za_data_7;
output 	za_data_6;
output 	za_data_20;
output 	za_data_19;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	sdram_wire_dq_0;
input 	sdram_wire_dq_1;
input 	sdram_wire_dq_2;
input 	sdram_wire_dq_3;
input 	sdram_wire_dq_4;
input 	sdram_wire_dq_5;
input 	sdram_wire_dq_6;
input 	sdram_wire_dq_7;
input 	sdram_wire_dq_8;
input 	sdram_wire_dq_9;
input 	sdram_wire_dq_10;
input 	sdram_wire_dq_11;
input 	sdram_wire_dq_12;
input 	sdram_wire_dq_13;
input 	sdram_wire_dq_14;
input 	sdram_wire_dq_15;
input 	sdram_wire_dq_16;
input 	sdram_wire_dq_17;
input 	sdram_wire_dq_18;
input 	sdram_wire_dq_19;
input 	sdram_wire_dq_20;
input 	sdram_wire_dq_21;
input 	sdram_wire_dq_22;
input 	sdram_wire_dq_23;
input 	sdram_wire_dq_24;
input 	sdram_wire_dq_25;
input 	sdram_wire_dq_26;
input 	sdram_wire_dq_27;
input 	sdram_wire_dq_28;
input 	sdram_wire_dq_29;
input 	sdram_wire_dq_30;
input 	sdram_wire_dq_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_address~q ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[56]~0_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[57]~1_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[58]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[58]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[59]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[59]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[46]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[46]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[60]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[60]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[47]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[47]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[48]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[48]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[49]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[49]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[61]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[61]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[50]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[50]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[51]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[51]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[52]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[52]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[53]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[53]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[54]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[54]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_1[55]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|entry_0[55]~q ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[36]~2_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[37]~3_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[38]~4_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[39]~5_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[40]~6_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[41]~7_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[42]~8_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[43]~9_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[44]~10_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[45]~11_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[46]~12_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[60]~13_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[32]~14_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[33]~15_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[34]~16_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[35]~17_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[47]~18_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[61]~19_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[58]~20_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[59]~21_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[48]~22_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[49]~23_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[50]~24_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[51]~25_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[52]~26_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[53]~27_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[54]~28_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[55]~29_combout ;
wire \comb~0_combout ;
wire \comb~1_combout ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[0]~30_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[1]~31_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[2]~32_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[3]~33_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[4]~34_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[5]~35_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[6]~36_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[7]~37_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[8]~38_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[9]~39_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[10]~40_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[11]~41_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[12]~42_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[13]~43_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[14]~44_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[15]~45_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[16]~46_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[17]~47_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[18]~48_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[19]~49_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[20]~50_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[21]~51_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[22]~52_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[23]~53_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[24]~54_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[25]~55_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[26]~56_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[27]~57_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[28]~58_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[29]~59_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[30]~60_combout ;
wire \the_sdram_demo_sdram_input_efifo_module|rd_data[31]~61_combout ;
wire \active_addr[20]~q ;
wire \active_addr[21]~q ;
wire \active_addr[22]~q ;
wire \Equal3~0_combout ;
wire \active_addr[23]~q ;
wire \Equal3~1_combout ;
wire \pending~0_combout ;
wire \active_addr[10]~q ;
wire \Equal2~0_combout ;
wire \active_addr[24]~q ;
wire \Equal2~1_combout ;
wire \active_addr[11]~q ;
wire \Equal3~2_combout ;
wire \active_addr[12]~q ;
wire \Equal3~3_combout ;
wire \active_addr[13]~q ;
wire \Equal3~4_combout ;
wire \active_rnw~q ;
wire \Add0~9_sumout ;
wire \refresh_counter~0_combout ;
wire \refresh_counter[0]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \refresh_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~49_sumout ;
wire \refresh_counter[2]~q ;
wire \Add0~50 ;
wire \Add0~45_sumout ;
wire \refresh_counter~8_combout ;
wire \refresh_counter[3]~q ;
wire \Add0~46 ;
wire \Add0~41_sumout ;
wire \refresh_counter~7_combout ;
wire \refresh_counter[4]~q ;
wire \Add0~42 ;
wire \Add0~37_sumout ;
wire \refresh_counter~6_combout ;
wire \refresh_counter[5]~q ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \refresh_counter~5_combout ;
wire \refresh_counter[6]~q ;
wire \Add0~34 ;
wire \Add0~1_sumout ;
wire \refresh_counter[7]~9_combout ;
wire \refresh_counter[7]~q ;
wire \Add0~2 ;
wire \Add0~29_sumout ;
wire \refresh_counter[8]~12_combout ;
wire \refresh_counter[8]~q ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \refresh_counter~4_combout ;
wire \refresh_counter[9]~q ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \refresh_counter~3_combout ;
wire \refresh_counter[10]~q ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \refresh_counter~2_combout ;
wire \refresh_counter[11]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \refresh_counter~1_combout ;
wire \refresh_counter[12]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \i_count[1]~0_combout ;
wire \i_count[0]~2_combout ;
wire \i_count[0]~q ;
wire \i_count[1]~1_combout ;
wire \i_count[1]~q ;
wire \WideOr6~combout ;
wire \i_next.000~0_combout ;
wire \i_next.000~q ;
wire \Selector7~0_combout ;
wire \i_state.000~q ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \i_count[2]~q ;
wire \Selector8~0_combout ;
wire \i_state.001~q ;
wire \Selector6~0_combout ;
wire \i_refs[0]~q ;
wire \Selector5~0_combout ;
wire \i_refs[1]~q ;
wire \Selector4~0_combout ;
wire \i_refs[2]~q ;
wire \Selector18~0_combout ;
wire \Selector16~0_combout ;
wire \i_next.010~q ;
wire \Selector9~0_combout ;
wire \i_state.010~q ;
wire \Selector18~1_combout ;
wire \i_next.111~q ;
wire \Selector12~0_combout ;
wire \i_state.111~q ;
wire \Selector10~0_combout ;
wire \i_state.011~q ;
wire \Selector17~0_combout ;
wire \i_next.101~q ;
wire \i_state.101~0_combout ;
wire \i_state.101~q ;
wire \init_done~0_combout ;
wire \init_done~q ;
wire \Selector32~0_combout ;
wire \m_state.100000000~q ;
wire \active_addr[14]~q ;
wire \Equal3~5_combout ;
wire \active_addr[15]~q ;
wire \Equal3~6_combout ;
wire \active_addr[16]~q ;
wire \Equal3~7_combout ;
wire \active_addr[17]~q ;
wire \Equal3~8_combout ;
wire \active_addr[18]~q ;
wire \Equal3~9_combout ;
wire \active_addr[19]~q ;
wire \Equal3~10_combout ;
wire \pending~3_combout ;
wire \pending~4_combout ;
wire \m_next~17_combout ;
wire \Selector35~0_combout ;
wire \Selector35~1_combout ;
wire \Selector34~0_combout ;
wire \Selector34~1_combout ;
wire \m_next.000001000~q ;
wire \Selector28~0_combout ;
wire \Selector28~1_combout ;
wire \Selector29~0_combout ;
wire \m_state.000100000~q ;
wire \Selector24~1_combout ;
wire \Selector30~1_combout ;
wire \m_state.001000000~q ;
wire \Selector36~2_combout ;
wire \Selector28~3_combout ;
wire \Selector28~4_combout ;
wire \Selector28~5_combout ;
wire \Selector35~2_combout ;
wire \Selector35~3_combout ;
wire \m_next.000010000~q ;
wire \Selector28~6_combout ;
wire \m_state.000010000~q ;
wire \Selector38~0_combout ;
wire \Selector38~1_combout ;
wire \Selector39~0_combout ;
wire \Selector39~1_combout ;
wire \Selector39~2_combout ;
wire \Selector39~3_combout ;
wire \Selector39~4_combout ;
wire \Selector39~5_combout ;
wire \m_count[0]~q ;
wire \Selector38~2_combout ;
wire \Selector38~3_combout ;
wire \Selector38~4_combout ;
wire \m_count[1]~q ;
wire \Selector24~0_combout ;
wire \Selector28~2_combout ;
wire \Selector27~0_combout ;
wire \m_state.000001000~q ;
wire \WideOr9~0_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \m_state.000000100~q ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \m_next.010000000~q ;
wire \Selector24~2_combout ;
wire \Selector24~3_combout ;
wire \Selector31~0_combout ;
wire \m_state.010000000~q ;
wire \Selector23~0_combout ;
wire \ack_refresh_request~q ;
wire \refresh_request~0_combout ;
wire \refresh_request~q ;
wire \Selector25~0_combout ;
wire \m_state.000000010~q ;
wire \WideOr8~0_combout ;
wire \Selector33~0_combout ;
wire \Selector33~1_combout ;
wire \Selector33~2_combout ;
wire \m_next.000000001~q ;
wire \Selector24~4_combout ;
wire \m_state.000000001~q ;
wire \Selector30~0_combout ;
wire \active_cs_n~0_combout ;
wire \active_cs_n~q ;
wire \pending~1_combout ;
wire \pending~2_combout ;
wire \Selector41~0_combout ;
wire \active_rnw~0_combout ;
wire \active_rnw~1_combout ;
wire \active_rnw~2_combout ;
wire \active_addr[0]~q ;
wire \Selector41~1_combout ;
wire \f_pop~q ;
wire \m_addr[6]~0_combout ;
wire \i_addr[12]~q ;
wire \Selector116~0_combout ;
wire \m_addr[6]~1_combout ;
wire \active_addr[1]~q ;
wire \Selector115~0_combout ;
wire \active_addr[2]~q ;
wire \Selector114~0_combout ;
wire \active_addr[3]~q ;
wire \Selector113~0_combout ;
wire \active_addr[6]~q ;
wire \Selector110~0_combout ;
wire \active_addr[7]~q ;
wire \Selector109~0_combout ;
wire \active_addr[8]~q ;
wire \Selector108~0_combout ;
wire \active_addr[9]~q ;
wire \Selector107~0_combout ;
wire \always5~0_combout ;
wire \active_addr[4]~q ;
wire \Selector112~0_combout ;
wire \Selector112~1_combout ;
wire \active_addr[5]~q ;
wire \Selector111~0_combout ;
wire \Selector106~0_combout ;
wire \Selector105~0_combout ;
wire \Selector104~0_combout ;
wire \Selector118~0_combout ;
wire \WideOr16~0_combout ;
wire \Selector117~0_combout ;
wire \Selector2~0_combout ;
wire \i_cmd[1]~q ;
wire \Selector21~0_combout ;
wire \Selector0~0_combout ;
wire \i_cmd[3]~q ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \active_dqm[0]~q ;
wire \Selector154~0_combout ;
wire \active_dqm[1]~q ;
wire \Selector153~0_combout ;
wire \active_dqm[2]~q ;
wire \Selector152~0_combout ;
wire \active_dqm[3]~q ;
wire \Selector151~0_combout ;
wire \Selector1~0_combout ;
wire \i_cmd[2]~q ;
wire \Selector20~0_combout ;
wire \Selector3~0_combout ;
wire \i_cmd[0]~q ;
wire \Selector22~0_combout ;
wire \Equal4~0_combout ;
wire \rd_valid[0]~q ;
wire \rd_valid[1]~q ;
wire \rd_valid[2]~q ;
wire \m_data[1]~0_combout ;
wire \active_data[0]~q ;
wire \WideOr17~0_combout ;
wire \Selector150~0_combout ;
wire \active_data[1]~q ;
wire \Selector149~0_combout ;
wire \active_data[2]~q ;
wire \Selector148~0_combout ;
wire \active_data[3]~q ;
wire \Selector147~0_combout ;
wire \active_data[4]~q ;
wire \Selector146~0_combout ;
wire \active_data[5]~q ;
wire \Selector145~0_combout ;
wire \active_data[6]~q ;
wire \Selector144~0_combout ;
wire \active_data[7]~q ;
wire \Selector143~0_combout ;
wire \active_data[8]~q ;
wire \Selector142~0_combout ;
wire \active_data[9]~q ;
wire \Selector141~0_combout ;
wire \active_data[10]~q ;
wire \Selector140~0_combout ;
wire \active_data[11]~q ;
wire \Selector139~0_combout ;
wire \active_data[12]~q ;
wire \Selector138~0_combout ;
wire \active_data[13]~q ;
wire \Selector137~0_combout ;
wire \active_data[14]~q ;
wire \Selector136~0_combout ;
wire \active_data[15]~q ;
wire \Selector135~0_combout ;
wire \active_data[16]~q ;
wire \Selector134~0_combout ;
wire \active_data[17]~q ;
wire \Selector133~0_combout ;
wire \active_data[18]~q ;
wire \Selector132~0_combout ;
wire \active_data[19]~q ;
wire \Selector131~0_combout ;
wire \active_data[20]~q ;
wire \Selector130~0_combout ;
wire \active_data[21]~q ;
wire \Selector129~0_combout ;
wire \active_data[22]~q ;
wire \Selector128~0_combout ;
wire \active_data[23]~q ;
wire \Selector127~0_combout ;
wire \active_data[24]~q ;
wire \Selector126~0_combout ;
wire \active_data[25]~q ;
wire \Selector125~0_combout ;
wire \active_data[26]~q ;
wire \Selector124~0_combout ;
wire \active_data[27]~q ;
wire \Selector123~0_combout ;
wire \active_data[28]~q ;
wire \Selector122~0_combout ;
wire \active_data[29]~q ;
wire \Selector121~0_combout ;
wire \active_data[30]~q ;
wire \Selector120~0_combout ;
wire \active_data[31]~q ;
wire \Selector119~0_combout ;


sdram_demo_sdram_demo_sdram_input_efifo_module the_sdram_demo_sdram_input_efifo_module(
	.reset_n(r_sync_rst),
	.always0(always0),
	.f_pop(\f_pop~q ),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.Equal1(\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.rd_address1(\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.rd_data_56(\the_sdram_demo_sdram_input_efifo_module|rd_data[56]~0_combout ),
	.rd_data_57(\the_sdram_demo_sdram_input_efifo_module|rd_data[57]~1_combout ),
	.entry_1_58(\the_sdram_demo_sdram_input_efifo_module|entry_1[58]~q ),
	.entry_0_58(\the_sdram_demo_sdram_input_efifo_module|entry_0[58]~q ),
	.entry_1_59(\the_sdram_demo_sdram_input_efifo_module|entry_1[59]~q ),
	.entry_0_59(\the_sdram_demo_sdram_input_efifo_module|entry_0[59]~q ),
	.entry_1_46(\the_sdram_demo_sdram_input_efifo_module|entry_1[46]~q ),
	.entry_0_46(\the_sdram_demo_sdram_input_efifo_module|entry_0[46]~q ),
	.entry_1_60(\the_sdram_demo_sdram_input_efifo_module|entry_1[60]~q ),
	.entry_0_60(\the_sdram_demo_sdram_input_efifo_module|entry_0[60]~q ),
	.entry_1_47(\the_sdram_demo_sdram_input_efifo_module|entry_1[47]~q ),
	.entry_0_47(\the_sdram_demo_sdram_input_efifo_module|entry_0[47]~q ),
	.entry_1_48(\the_sdram_demo_sdram_input_efifo_module|entry_1[48]~q ),
	.entry_0_48(\the_sdram_demo_sdram_input_efifo_module|entry_0[48]~q ),
	.entry_1_49(\the_sdram_demo_sdram_input_efifo_module|entry_1[49]~q ),
	.entry_0_49(\the_sdram_demo_sdram_input_efifo_module|entry_0[49]~q ),
	.entry_1_61(\the_sdram_demo_sdram_input_efifo_module|entry_1[61]~q ),
	.entry_0_61(\the_sdram_demo_sdram_input_efifo_module|entry_0[61]~q ),
	.entry_1_50(\the_sdram_demo_sdram_input_efifo_module|entry_1[50]~q ),
	.entry_0_50(\the_sdram_demo_sdram_input_efifo_module|entry_0[50]~q ),
	.entry_1_51(\the_sdram_demo_sdram_input_efifo_module|entry_1[51]~q ),
	.entry_0_51(\the_sdram_demo_sdram_input_efifo_module|entry_0[51]~q ),
	.entry_1_52(\the_sdram_demo_sdram_input_efifo_module|entry_1[52]~q ),
	.entry_0_52(\the_sdram_demo_sdram_input_efifo_module|entry_0[52]~q ),
	.entry_1_53(\the_sdram_demo_sdram_input_efifo_module|entry_1[53]~q ),
	.entry_0_53(\the_sdram_demo_sdram_input_efifo_module|entry_0[53]~q ),
	.entry_1_54(\the_sdram_demo_sdram_input_efifo_module|entry_1[54]~q ),
	.entry_0_54(\the_sdram_demo_sdram_input_efifo_module|entry_0[54]~q ),
	.entry_1_55(\the_sdram_demo_sdram_input_efifo_module|entry_1[55]~q ),
	.entry_0_55(\the_sdram_demo_sdram_input_efifo_module|entry_0[55]~q ),
	.Selector41(\Selector41~0_combout ),
	.rd_data_36(\the_sdram_demo_sdram_input_efifo_module|rd_data[36]~2_combout ),
	.rd_data_37(\the_sdram_demo_sdram_input_efifo_module|rd_data[37]~3_combout ),
	.rd_data_38(\the_sdram_demo_sdram_input_efifo_module|rd_data[38]~4_combout ),
	.rd_data_39(\the_sdram_demo_sdram_input_efifo_module|rd_data[39]~5_combout ),
	.rd_data_40(\the_sdram_demo_sdram_input_efifo_module|rd_data[40]~6_combout ),
	.rd_data_41(\the_sdram_demo_sdram_input_efifo_module|rd_data[41]~7_combout ),
	.rd_data_42(\the_sdram_demo_sdram_input_efifo_module|rd_data[42]~8_combout ),
	.rd_data_43(\the_sdram_demo_sdram_input_efifo_module|rd_data[43]~9_combout ),
	.rd_data_44(\the_sdram_demo_sdram_input_efifo_module|rd_data[44]~10_combout ),
	.rd_data_45(\the_sdram_demo_sdram_input_efifo_module|rd_data[45]~11_combout ),
	.rd_data_46(\the_sdram_demo_sdram_input_efifo_module|rd_data[46]~12_combout ),
	.rd_data_60(\the_sdram_demo_sdram_input_efifo_module|rd_data[60]~13_combout ),
	.rd_data_32(\the_sdram_demo_sdram_input_efifo_module|rd_data[32]~14_combout ),
	.rd_data_33(\the_sdram_demo_sdram_input_efifo_module|rd_data[33]~15_combout ),
	.rd_data_34(\the_sdram_demo_sdram_input_efifo_module|rd_data[34]~16_combout ),
	.rd_data_35(\the_sdram_demo_sdram_input_efifo_module|rd_data[35]~17_combout ),
	.saved_grant_0(saved_grant_0),
	.WideOr0(WideOr0),
	.rd_data_47(\the_sdram_demo_sdram_input_efifo_module|rd_data[47]~18_combout ),
	.rd_data_61(\the_sdram_demo_sdram_input_efifo_module|rd_data[61]~19_combout ),
	.Equal11(Equal1),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.src_data_68(src_data_68),
	.src_data_58(src_data_58),
	.src_valid1(src_valid1),
	.src_data_59(src_data_59),
	.rd_data_58(\the_sdram_demo_sdram_input_efifo_module|rd_data[58]~20_combout ),
	.src_data_60(src_data_60),
	.rd_data_59(\the_sdram_demo_sdram_input_efifo_module|rd_data[59]~21_combout ),
	.src_data_61(src_data_61),
	.src_data_48(src_data_48),
	.src_data_62(src_data_62),
	.src_data_49(src_data_49),
	.rd_data_48(\the_sdram_demo_sdram_input_efifo_module|rd_data[48]~22_combout ),
	.src_data_50(src_data_50),
	.rd_data_49(\the_sdram_demo_sdram_input_efifo_module|rd_data[49]~23_combout ),
	.src_data_51(src_data_51),
	.m0_write(m0_write1),
	.rd_data_50(\the_sdram_demo_sdram_input_efifo_module|rd_data[50]~24_combout ),
	.src_data_52(src_data_52),
	.rd_data_51(\the_sdram_demo_sdram_input_efifo_module|rd_data[51]~25_combout ),
	.src_data_53(src_data_53),
	.rd_data_52(\the_sdram_demo_sdram_input_efifo_module|rd_data[52]~26_combout ),
	.src_data_54(src_data_54),
	.rd_data_53(\the_sdram_demo_sdram_input_efifo_module|rd_data[53]~27_combout ),
	.src_data_55(src_data_55),
	.rd_data_54(\the_sdram_demo_sdram_input_efifo_module|rd_data[54]~28_combout ),
	.src_data_56(src_data_56),
	.rd_data_55(\the_sdram_demo_sdram_input_efifo_module|rd_data[55]~29_combout ),
	.src_data_57(src_data_57),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.comb(\comb~0_combout ),
	.comb1(\comb~1_combout ),
	.comb2(\comb~2_combout ),
	.comb3(\comb~3_combout ),
	.rd_data_0(\the_sdram_demo_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.rd_data_1(\the_sdram_demo_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.rd_data_2(\the_sdram_demo_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.rd_data_3(\the_sdram_demo_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.rd_data_4(\the_sdram_demo_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.rd_data_5(\the_sdram_demo_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.rd_data_6(\the_sdram_demo_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.rd_data_7(\the_sdram_demo_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.rd_data_8(\the_sdram_demo_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.rd_data_9(\the_sdram_demo_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.rd_data_10(\the_sdram_demo_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.rd_data_11(\the_sdram_demo_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.rd_data_12(\the_sdram_demo_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.rd_data_13(\the_sdram_demo_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.rd_data_14(\the_sdram_demo_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.rd_data_15(\the_sdram_demo_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.rd_data_16(\the_sdram_demo_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.rd_data_17(\the_sdram_demo_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.rd_data_18(\the_sdram_demo_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.rd_data_19(\the_sdram_demo_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.rd_data_20(\the_sdram_demo_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.rd_data_21(\the_sdram_demo_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.rd_data_22(\the_sdram_demo_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.rd_data_23(\the_sdram_demo_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.rd_data_24(\the_sdram_demo_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.rd_data_25(\the_sdram_demo_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.rd_data_26(\the_sdram_demo_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.rd_data_27(\the_sdram_demo_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.rd_data_28(\the_sdram_demo_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.rd_data_29(\the_sdram_demo_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.rd_data_30(\the_sdram_demo_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.rd_data_31(\the_sdram_demo_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.clk(clk_clk));

cyclonev_lcell_comb \comb~0 (
	.dataa(!src_valid1),
	.datab(!saved_grant_1),
	.datac(!src_valid),
	.datad(!d_byteenable_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~1 (
	.dataa(!src_valid1),
	.datab(!saved_grant_1),
	.datac(!src_valid),
	.datad(!m0_write),
	.datae(!d_byteenable_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~1 .extended_lut = "off";
defparam \comb~1 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \comb~1 .shared_arith = "off";

cyclonev_lcell_comb \comb~2 (
	.dataa(!src_valid1),
	.datab(!saved_grant_1),
	.datac(!src_valid),
	.datad(!m0_write),
	.datae(!d_byteenable_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~2 .extended_lut = "off";
defparam \comb~2 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \comb~2 .shared_arith = "off";

cyclonev_lcell_comb \comb~3 (
	.dataa(!src_valid1),
	.datab(!saved_grant_1),
	.datac(!src_valid),
	.datad(!m0_write),
	.datae(!d_byteenable_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~3 .extended_lut = "off";
defparam \comb~3 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \comb~3 .shared_arith = "off";

dffeas \m_addr[0] (
	.clk(clk_clk),
	.d(\Selector116~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_0),
	.prn(vcc));
defparam \m_addr[0] .is_wysiwyg = "true";
defparam \m_addr[0] .power_up = "low";

dffeas \m_addr[1] (
	.clk(clk_clk),
	.d(\Selector115~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_1),
	.prn(vcc));
defparam \m_addr[1] .is_wysiwyg = "true";
defparam \m_addr[1] .power_up = "low";

dffeas \m_addr[2] (
	.clk(clk_clk),
	.d(\Selector114~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_2),
	.prn(vcc));
defparam \m_addr[2] .is_wysiwyg = "true";
defparam \m_addr[2] .power_up = "low";

dffeas \m_addr[3] (
	.clk(clk_clk),
	.d(\Selector113~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_3),
	.prn(vcc));
defparam \m_addr[3] .is_wysiwyg = "true";
defparam \m_addr[3] .power_up = "low";

dffeas \m_addr[6] (
	.clk(clk_clk),
	.d(\Selector110~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_6),
	.prn(vcc));
defparam \m_addr[6] .is_wysiwyg = "true";
defparam \m_addr[6] .power_up = "low";

dffeas \m_addr[7] (
	.clk(clk_clk),
	.d(\Selector109~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_7),
	.prn(vcc));
defparam \m_addr[7] .is_wysiwyg = "true";
defparam \m_addr[7] .power_up = "low";

dffeas \m_addr[8] (
	.clk(clk_clk),
	.d(\Selector108~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_8),
	.prn(vcc));
defparam \m_addr[8] .is_wysiwyg = "true";
defparam \m_addr[8] .power_up = "low";

dffeas \m_addr[9] (
	.clk(clk_clk),
	.d(\Selector107~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_9),
	.prn(vcc));
defparam \m_addr[9] .is_wysiwyg = "true";
defparam \m_addr[9] .power_up = "low";

dffeas oe(
	.clk(clk_clk),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\m_state.000010000~q ),
	.sload(gnd),
	.ena(vcc),
	.q(oe1),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

dffeas \m_addr[4] (
	.clk(clk_clk),
	.d(\Selector112~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_4),
	.prn(vcc));
defparam \m_addr[4] .is_wysiwyg = "true";
defparam \m_addr[4] .power_up = "low";

dffeas \m_addr[5] (
	.clk(clk_clk),
	.d(\Selector111~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_5),
	.prn(vcc));
defparam \m_addr[5] .is_wysiwyg = "true";
defparam \m_addr[5] .power_up = "low";

dffeas \m_addr[10] (
	.clk(clk_clk),
	.d(\Selector106~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_10),
	.prn(vcc));
defparam \m_addr[10] .is_wysiwyg = "true";
defparam \m_addr[10] .power_up = "low";

dffeas \m_addr[11] (
	.clk(clk_clk),
	.d(\Selector105~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_11),
	.prn(vcc));
defparam \m_addr[11] .is_wysiwyg = "true";
defparam \m_addr[11] .power_up = "low";

dffeas \m_addr[12] (
	.clk(clk_clk),
	.d(\Selector104~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[6]~1_combout ),
	.q(m_addr_12),
	.prn(vcc));
defparam \m_addr[12] .is_wysiwyg = "true";
defparam \m_addr[12] .power_up = "low";

dffeas \m_bank[0] (
	.clk(clk_clk),
	.d(\Selector118~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_0),
	.prn(vcc));
defparam \m_bank[0] .is_wysiwyg = "true";
defparam \m_bank[0] .power_up = "low";

dffeas \m_bank[1] (
	.clk(clk_clk),
	.d(\Selector117~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_1),
	.prn(vcc));
defparam \m_bank[1] .is_wysiwyg = "true";
defparam \m_bank[1] .power_up = "low";

dffeas \m_cmd[1] (
	.clk(clk_clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_1),
	.prn(vcc));
defparam \m_cmd[1] .is_wysiwyg = "true";
defparam \m_cmd[1] .power_up = "low";

dffeas \m_cmd[3] (
	.clk(clk_clk),
	.d(\Selector19~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_3),
	.prn(vcc));
defparam \m_cmd[3] .is_wysiwyg = "true";
defparam \m_cmd[3] .power_up = "low";

dffeas \m_dqm[0] (
	.clk(clk_clk),
	.d(\Selector154~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_0),
	.prn(vcc));
defparam \m_dqm[0] .is_wysiwyg = "true";
defparam \m_dqm[0] .power_up = "low";

dffeas \m_dqm[1] (
	.clk(clk_clk),
	.d(\Selector153~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_1),
	.prn(vcc));
defparam \m_dqm[1] .is_wysiwyg = "true";
defparam \m_dqm[1] .power_up = "low";

dffeas \m_dqm[2] (
	.clk(clk_clk),
	.d(\Selector152~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_2),
	.prn(vcc));
defparam \m_dqm[2] .is_wysiwyg = "true";
defparam \m_dqm[2] .power_up = "low";

dffeas \m_dqm[3] (
	.clk(clk_clk),
	.d(\Selector151~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_3),
	.prn(vcc));
defparam \m_dqm[3] .is_wysiwyg = "true";
defparam \m_dqm[3] .power_up = "low";

dffeas \m_cmd[2] (
	.clk(clk_clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_2),
	.prn(vcc));
defparam \m_cmd[2] .is_wysiwyg = "true";
defparam \m_cmd[2] .power_up = "low";

dffeas \m_cmd[0] (
	.clk(clk_clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_0),
	.prn(vcc));
defparam \m_cmd[0] .is_wysiwyg = "true";
defparam \m_cmd[0] .power_up = "low";

dffeas za_valid(
	.clk(clk_clk),
	.d(\rd_valid[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_valid1),
	.prn(vcc));
defparam za_valid.is_wysiwyg = "true";
defparam za_valid.power_up = "low";

dffeas \m_data[0] (
	.clk(clk_clk),
	.d(\Selector150~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_0),
	.prn(vcc));
defparam \m_data[0] .is_wysiwyg = "true";
defparam \m_data[0] .power_up = "low";

dffeas \m_data[1] (
	.clk(clk_clk),
	.d(\Selector149~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_1),
	.prn(vcc));
defparam \m_data[1] .is_wysiwyg = "true";
defparam \m_data[1] .power_up = "low";

dffeas \m_data[2] (
	.clk(clk_clk),
	.d(\Selector148~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_2),
	.prn(vcc));
defparam \m_data[2] .is_wysiwyg = "true";
defparam \m_data[2] .power_up = "low";

dffeas \m_data[3] (
	.clk(clk_clk),
	.d(\Selector147~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_3),
	.prn(vcc));
defparam \m_data[3] .is_wysiwyg = "true";
defparam \m_data[3] .power_up = "low";

dffeas \m_data[4] (
	.clk(clk_clk),
	.d(\Selector146~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_4),
	.prn(vcc));
defparam \m_data[4] .is_wysiwyg = "true";
defparam \m_data[4] .power_up = "low";

dffeas \m_data[5] (
	.clk(clk_clk),
	.d(\Selector145~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_5),
	.prn(vcc));
defparam \m_data[5] .is_wysiwyg = "true";
defparam \m_data[5] .power_up = "low";

dffeas \m_data[6] (
	.clk(clk_clk),
	.d(\Selector144~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_6),
	.prn(vcc));
defparam \m_data[6] .is_wysiwyg = "true";
defparam \m_data[6] .power_up = "low";

dffeas \m_data[7] (
	.clk(clk_clk),
	.d(\Selector143~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_7),
	.prn(vcc));
defparam \m_data[7] .is_wysiwyg = "true";
defparam \m_data[7] .power_up = "low";

dffeas \m_data[8] (
	.clk(clk_clk),
	.d(\Selector142~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_8),
	.prn(vcc));
defparam \m_data[8] .is_wysiwyg = "true";
defparam \m_data[8] .power_up = "low";

dffeas \m_data[9] (
	.clk(clk_clk),
	.d(\Selector141~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_9),
	.prn(vcc));
defparam \m_data[9] .is_wysiwyg = "true";
defparam \m_data[9] .power_up = "low";

dffeas \m_data[10] (
	.clk(clk_clk),
	.d(\Selector140~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_10),
	.prn(vcc));
defparam \m_data[10] .is_wysiwyg = "true";
defparam \m_data[10] .power_up = "low";

dffeas \m_data[11] (
	.clk(clk_clk),
	.d(\Selector139~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_11),
	.prn(vcc));
defparam \m_data[11] .is_wysiwyg = "true";
defparam \m_data[11] .power_up = "low";

dffeas \m_data[12] (
	.clk(clk_clk),
	.d(\Selector138~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_12),
	.prn(vcc));
defparam \m_data[12] .is_wysiwyg = "true";
defparam \m_data[12] .power_up = "low";

dffeas \m_data[13] (
	.clk(clk_clk),
	.d(\Selector137~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_13),
	.prn(vcc));
defparam \m_data[13] .is_wysiwyg = "true";
defparam \m_data[13] .power_up = "low";

dffeas \m_data[14] (
	.clk(clk_clk),
	.d(\Selector136~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_14),
	.prn(vcc));
defparam \m_data[14] .is_wysiwyg = "true";
defparam \m_data[14] .power_up = "low";

dffeas \m_data[15] (
	.clk(clk_clk),
	.d(\Selector135~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_15),
	.prn(vcc));
defparam \m_data[15] .is_wysiwyg = "true";
defparam \m_data[15] .power_up = "low";

dffeas \m_data[16] (
	.clk(clk_clk),
	.d(\Selector134~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_16),
	.prn(vcc));
defparam \m_data[16] .is_wysiwyg = "true";
defparam \m_data[16] .power_up = "low";

dffeas \m_data[17] (
	.clk(clk_clk),
	.d(\Selector133~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_17),
	.prn(vcc));
defparam \m_data[17] .is_wysiwyg = "true";
defparam \m_data[17] .power_up = "low";

dffeas \m_data[18] (
	.clk(clk_clk),
	.d(\Selector132~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_18),
	.prn(vcc));
defparam \m_data[18] .is_wysiwyg = "true";
defparam \m_data[18] .power_up = "low";

dffeas \m_data[19] (
	.clk(clk_clk),
	.d(\Selector131~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_19),
	.prn(vcc));
defparam \m_data[19] .is_wysiwyg = "true";
defparam \m_data[19] .power_up = "low";

dffeas \m_data[20] (
	.clk(clk_clk),
	.d(\Selector130~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_20),
	.prn(vcc));
defparam \m_data[20] .is_wysiwyg = "true";
defparam \m_data[20] .power_up = "low";

dffeas \m_data[21] (
	.clk(clk_clk),
	.d(\Selector129~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_21),
	.prn(vcc));
defparam \m_data[21] .is_wysiwyg = "true";
defparam \m_data[21] .power_up = "low";

dffeas \m_data[22] (
	.clk(clk_clk),
	.d(\Selector128~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_22),
	.prn(vcc));
defparam \m_data[22] .is_wysiwyg = "true";
defparam \m_data[22] .power_up = "low";

dffeas \m_data[23] (
	.clk(clk_clk),
	.d(\Selector127~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_23),
	.prn(vcc));
defparam \m_data[23] .is_wysiwyg = "true";
defparam \m_data[23] .power_up = "low";

dffeas \m_data[24] (
	.clk(clk_clk),
	.d(\Selector126~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_24),
	.prn(vcc));
defparam \m_data[24] .is_wysiwyg = "true";
defparam \m_data[24] .power_up = "low";

dffeas \m_data[25] (
	.clk(clk_clk),
	.d(\Selector125~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_25),
	.prn(vcc));
defparam \m_data[25] .is_wysiwyg = "true";
defparam \m_data[25] .power_up = "low";

dffeas \m_data[26] (
	.clk(clk_clk),
	.d(\Selector124~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_26),
	.prn(vcc));
defparam \m_data[26] .is_wysiwyg = "true";
defparam \m_data[26] .power_up = "low";

dffeas \m_data[27] (
	.clk(clk_clk),
	.d(\Selector123~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_27),
	.prn(vcc));
defparam \m_data[27] .is_wysiwyg = "true";
defparam \m_data[27] .power_up = "low";

dffeas \m_data[28] (
	.clk(clk_clk),
	.d(\Selector122~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_28),
	.prn(vcc));
defparam \m_data[28] .is_wysiwyg = "true";
defparam \m_data[28] .power_up = "low";

dffeas \m_data[29] (
	.clk(clk_clk),
	.d(\Selector121~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_29),
	.prn(vcc));
defparam \m_data[29] .is_wysiwyg = "true";
defparam \m_data[29] .power_up = "low";

dffeas \m_data[30] (
	.clk(clk_clk),
	.d(\Selector120~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_30),
	.prn(vcc));
defparam \m_data[30] .is_wysiwyg = "true";
defparam \m_data[30] .power_up = "low";

dffeas \m_data[31] (
	.clk(clk_clk),
	.d(\Selector119~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_31),
	.prn(vcc));
defparam \m_data[31] .is_wysiwyg = "true";
defparam \m_data[31] .power_up = "low";

dffeas \za_data[0] (
	.clk(clk_clk),
	.d(sdram_wire_dq_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_0),
	.prn(vcc));
defparam \za_data[0] .is_wysiwyg = "true";
defparam \za_data[0] .power_up = "low";

dffeas \za_data[22] (
	.clk(clk_clk),
	.d(sdram_wire_dq_22),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_22),
	.prn(vcc));
defparam \za_data[22] .is_wysiwyg = "true";
defparam \za_data[22] .power_up = "low";

dffeas \za_data[23] (
	.clk(clk_clk),
	.d(sdram_wire_dq_23),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_23),
	.prn(vcc));
defparam \za_data[23] .is_wysiwyg = "true";
defparam \za_data[23] .power_up = "low";

dffeas \za_data[24] (
	.clk(clk_clk),
	.d(sdram_wire_dq_24),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_24),
	.prn(vcc));
defparam \za_data[24] .is_wysiwyg = "true";
defparam \za_data[24] .power_up = "low";

dffeas \za_data[25] (
	.clk(clk_clk),
	.d(sdram_wire_dq_25),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_25),
	.prn(vcc));
defparam \za_data[25] .is_wysiwyg = "true";
defparam \za_data[25] .power_up = "low";

dffeas \za_data[26] (
	.clk(clk_clk),
	.d(sdram_wire_dq_26),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_26),
	.prn(vcc));
defparam \za_data[26] .is_wysiwyg = "true";
defparam \za_data[26] .power_up = "low";

dffeas \za_data[1] (
	.clk(clk_clk),
	.d(sdram_wire_dq_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_1),
	.prn(vcc));
defparam \za_data[1] .is_wysiwyg = "true";
defparam \za_data[1] .power_up = "low";

dffeas \za_data[4] (
	.clk(clk_clk),
	.d(sdram_wire_dq_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_4),
	.prn(vcc));
defparam \za_data[4] .is_wysiwyg = "true";
defparam \za_data[4] .power_up = "low";

dffeas \za_data[3] (
	.clk(clk_clk),
	.d(sdram_wire_dq_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_3),
	.prn(vcc));
defparam \za_data[3] .is_wysiwyg = "true";
defparam \za_data[3] .power_up = "low";

dffeas \za_data[2] (
	.clk(clk_clk),
	.d(sdram_wire_dq_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_2),
	.prn(vcc));
defparam \za_data[2] .is_wysiwyg = "true";
defparam \za_data[2] .power_up = "low";

dffeas \za_data[11] (
	.clk(clk_clk),
	.d(sdram_wire_dq_11),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_11),
	.prn(vcc));
defparam \za_data[11] .is_wysiwyg = "true";
defparam \za_data[11] .power_up = "low";

dffeas \za_data[12] (
	.clk(clk_clk),
	.d(sdram_wire_dq_12),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_12),
	.prn(vcc));
defparam \za_data[12] .is_wysiwyg = "true";
defparam \za_data[12] .power_up = "low";

dffeas \za_data[13] (
	.clk(clk_clk),
	.d(sdram_wire_dq_13),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_13),
	.prn(vcc));
defparam \za_data[13] .is_wysiwyg = "true";
defparam \za_data[13] .power_up = "low";

dffeas \za_data[14] (
	.clk(clk_clk),
	.d(sdram_wire_dq_14),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_14),
	.prn(vcc));
defparam \za_data[14] .is_wysiwyg = "true";
defparam \za_data[14] .power_up = "low";

dffeas \za_data[15] (
	.clk(clk_clk),
	.d(sdram_wire_dq_15),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_15),
	.prn(vcc));
defparam \za_data[15] .is_wysiwyg = "true";
defparam \za_data[15] .power_up = "low";

dffeas \za_data[16] (
	.clk(clk_clk),
	.d(sdram_wire_dq_16),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_16),
	.prn(vcc));
defparam \za_data[16] .is_wysiwyg = "true";
defparam \za_data[16] .power_up = "low";

dffeas \za_data[5] (
	.clk(clk_clk),
	.d(sdram_wire_dq_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_5),
	.prn(vcc));
defparam \za_data[5] .is_wysiwyg = "true";
defparam \za_data[5] .power_up = "low";

dffeas \za_data[8] (
	.clk(clk_clk),
	.d(sdram_wire_dq_8),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_8),
	.prn(vcc));
defparam \za_data[8] .is_wysiwyg = "true";
defparam \za_data[8] .power_up = "low";

dffeas \za_data[10] (
	.clk(clk_clk),
	.d(sdram_wire_dq_10),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_10),
	.prn(vcc));
defparam \za_data[10] .is_wysiwyg = "true";
defparam \za_data[10] .power_up = "low";

dffeas \za_data[9] (
	.clk(clk_clk),
	.d(sdram_wire_dq_9),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_9),
	.prn(vcc));
defparam \za_data[9] .is_wysiwyg = "true";
defparam \za_data[9] .power_up = "low";

dffeas \za_data[28] (
	.clk(clk_clk),
	.d(sdram_wire_dq_28),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_28),
	.prn(vcc));
defparam \za_data[28] .is_wysiwyg = "true";
defparam \za_data[28] .power_up = "low";

dffeas \za_data[21] (
	.clk(clk_clk),
	.d(sdram_wire_dq_21),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_21),
	.prn(vcc));
defparam \za_data[21] .is_wysiwyg = "true";
defparam \za_data[21] .power_up = "low";

dffeas \za_data[29] (
	.clk(clk_clk),
	.d(sdram_wire_dq_29),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_29),
	.prn(vcc));
defparam \za_data[29] .is_wysiwyg = "true";
defparam \za_data[29] .power_up = "low";

dffeas \za_data[30] (
	.clk(clk_clk),
	.d(sdram_wire_dq_30),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_30),
	.prn(vcc));
defparam \za_data[30] .is_wysiwyg = "true";
defparam \za_data[30] .power_up = "low";

dffeas \za_data[31] (
	.clk(clk_clk),
	.d(sdram_wire_dq_31),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_31),
	.prn(vcc));
defparam \za_data[31] .is_wysiwyg = "true";
defparam \za_data[31] .power_up = "low";

dffeas \za_data[17] (
	.clk(clk_clk),
	.d(sdram_wire_dq_17),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_17),
	.prn(vcc));
defparam \za_data[17] .is_wysiwyg = "true";
defparam \za_data[17] .power_up = "low";

dffeas \za_data[18] (
	.clk(clk_clk),
	.d(sdram_wire_dq_18),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_18),
	.prn(vcc));
defparam \za_data[18] .is_wysiwyg = "true";
defparam \za_data[18] .power_up = "low";

dffeas \za_data[27] (
	.clk(clk_clk),
	.d(sdram_wire_dq_27),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_27),
	.prn(vcc));
defparam \za_data[27] .is_wysiwyg = "true";
defparam \za_data[27] .power_up = "low";

dffeas \za_data[7] (
	.clk(clk_clk),
	.d(sdram_wire_dq_7),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_7),
	.prn(vcc));
defparam \za_data[7] .is_wysiwyg = "true";
defparam \za_data[7] .power_up = "low";

dffeas \za_data[6] (
	.clk(clk_clk),
	.d(sdram_wire_dq_6),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_6),
	.prn(vcc));
defparam \za_data[6] .is_wysiwyg = "true";
defparam \za_data[6] .power_up = "low";

dffeas \za_data[20] (
	.clk(clk_clk),
	.d(sdram_wire_dq_20),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_20),
	.prn(vcc));
defparam \za_data[20] .is_wysiwyg = "true";
defparam \za_data[20] .power_up = "low";

dffeas \za_data[19] (
	.clk(clk_clk),
	.d(sdram_wire_dq_19),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_19),
	.prn(vcc));
defparam \za_data[19] .is_wysiwyg = "true";
defparam \za_data[19] .power_up = "low";

dffeas \active_addr[20] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[56]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[20]~q ),
	.prn(vcc));
defparam \active_addr[20] .is_wysiwyg = "true";
defparam \active_addr[20] .power_up = "low";

dffeas \active_addr[21] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[57]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[21]~q ),
	.prn(vcc));
defparam \active_addr[21] .is_wysiwyg = "true";
defparam \active_addr[21] .power_up = "low";

dffeas \active_addr[22] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[58]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[22]~q ),
	.prn(vcc));
defparam \active_addr[22] .is_wysiwyg = "true";
defparam \active_addr[22] .power_up = "low";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[22]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[58]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[58]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h6996699669966996;
defparam \Equal3~0 .shared_arith = "off";

dffeas \active_addr[23] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[59]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[23]~q ),
	.prn(vcc));
defparam \active_addr[23] .is_wysiwyg = "true";
defparam \active_addr[23] .power_up = "low";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[23]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[59]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[59]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'h6996699669966996;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \pending~0 (
	.dataa(!\active_addr[20]~q ),
	.datab(!\the_sdram_demo_sdram_input_efifo_module|rd_data[56]~0_combout ),
	.datac(!\active_addr[21]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[57]~1_combout ),
	.datae(!\Equal3~0_combout ),
	.dataf(!\Equal3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending~0 .extended_lut = "off";
defparam \pending~0 .lut_mask = 64'hFFFFFFFFFFFF6996;
defparam \pending~0 .shared_arith = "off";

dffeas \active_addr[10] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[46]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[10]~q ),
	.prn(vcc));
defparam \active_addr[10] .is_wysiwyg = "true";
defparam \active_addr[10] .power_up = "low";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[10]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[46]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[46]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h6996699669966996;
defparam \Equal2~0 .shared_arith = "off";

dffeas \active_addr[24] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[60]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[24]~q ),
	.prn(vcc));
defparam \active_addr[24] .is_wysiwyg = "true";
defparam \active_addr[24] .power_up = "low";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[24]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[60]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[60]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h6996699669966996;
defparam \Equal2~1 .shared_arith = "off";

dffeas \active_addr[11] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[47]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[11]~q ),
	.prn(vcc));
defparam \active_addr[11] .is_wysiwyg = "true";
defparam \active_addr[11] .power_up = "low";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[11]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[47]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[47]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'h6996699669966996;
defparam \Equal3~2 .shared_arith = "off";

dffeas \active_addr[12] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[48]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[12]~q ),
	.prn(vcc));
defparam \active_addr[12] .is_wysiwyg = "true";
defparam \active_addr[12] .power_up = "low";

cyclonev_lcell_comb \Equal3~3 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[12]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[48]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[48]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~3 .extended_lut = "off";
defparam \Equal3~3 .lut_mask = 64'h6996699669966996;
defparam \Equal3~3 .shared_arith = "off";

dffeas \active_addr[13] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[49]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[13]~q ),
	.prn(vcc));
defparam \active_addr[13] .is_wysiwyg = "true";
defparam \active_addr[13] .power_up = "low";

cyclonev_lcell_comb \Equal3~4 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[13]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[49]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[49]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~4 .extended_lut = "off";
defparam \Equal3~4 .lut_mask = 64'h6996699669966996;
defparam \Equal3~4 .shared_arith = "off";

dffeas active_rnw(
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[61]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_rnw~q ),
	.prn(vcc));
defparam active_rnw.is_wysiwyg = "true";
defparam active_rnw.power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~0 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~0 .extended_lut = "off";
defparam \refresh_counter~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~0 .shared_arith = "off";

dffeas \refresh_counter[0] (
	.clk(clk_clk),
	.d(\refresh_counter~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[0]~q ),
	.prn(vcc));
defparam \refresh_counter[0] .is_wysiwyg = "true";
defparam \refresh_counter[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \refresh_counter[1] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[1]~q ),
	.prn(vcc));
defparam \refresh_counter[1] .is_wysiwyg = "true";
defparam \refresh_counter[1] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \refresh_counter[2] (
	.clk(clk_clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[2]~q ),
	.prn(vcc));
defparam \refresh_counter[2] .is_wysiwyg = "true";
defparam \refresh_counter[2] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000000000FF00;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~8 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~8 .extended_lut = "off";
defparam \refresh_counter~8 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \refresh_counter~8 .shared_arith = "off";

dffeas \refresh_counter[3] (
	.clk(clk_clk),
	.d(\refresh_counter~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[3]~q ),
	.prn(vcc));
defparam \refresh_counter[3] .is_wysiwyg = "true";
defparam \refresh_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~7 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~41_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~7 .extended_lut = "off";
defparam \refresh_counter~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~7 .shared_arith = "off";

dffeas \refresh_counter[4] (
	.clk(clk_clk),
	.d(\refresh_counter~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[4]~q ),
	.prn(vcc));
defparam \refresh_counter[4] .is_wysiwyg = "true";
defparam \refresh_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~6 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~37_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~6 .extended_lut = "off";
defparam \refresh_counter~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~6 .shared_arith = "off";

dffeas \refresh_counter[5] (
	.clk(clk_clk),
	.d(\refresh_counter~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[5]~q ),
	.prn(vcc));
defparam \refresh_counter[5] .is_wysiwyg = "true";
defparam \refresh_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~5 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~33_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~5 .extended_lut = "off";
defparam \refresh_counter~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~5 .shared_arith = "off";

dffeas \refresh_counter[6] (
	.clk(clk_clk),
	.d(\refresh_counter~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[6]~q ),
	.prn(vcc));
defparam \refresh_counter[6] .is_wysiwyg = "true";
defparam \refresh_counter[6] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter[7]~9 (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter[7]~9 .extended_lut = "off";
defparam \refresh_counter[7]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \refresh_counter[7]~9 .shared_arith = "off";

dffeas \refresh_counter[7] (
	.clk(clk_clk),
	.d(\refresh_counter[7]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[7]~q ),
	.prn(vcc));
defparam \refresh_counter[7] .is_wysiwyg = "true";
defparam \refresh_counter[7] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000000000FF00;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter[8]~12 (
	.dataa(!\Add0~29_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter[8]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter[8]~12 .extended_lut = "off";
defparam \refresh_counter[8]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \refresh_counter[8]~12 .shared_arith = "off";

dffeas \refresh_counter[8] (
	.clk(clk_clk),
	.d(\refresh_counter[8]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[8]~q ),
	.prn(vcc));
defparam \refresh_counter[8] .is_wysiwyg = "true";
defparam \refresh_counter[8] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~4 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~25_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~4 .extended_lut = "off";
defparam \refresh_counter~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \refresh_counter~4 .shared_arith = "off";

dffeas \refresh_counter[9] (
	.clk(clk_clk),
	.d(\refresh_counter~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[9]~q ),
	.prn(vcc));
defparam \refresh_counter[9] .is_wysiwyg = "true";
defparam \refresh_counter[9] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~3 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~3 .extended_lut = "off";
defparam \refresh_counter~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~3 .shared_arith = "off";

dffeas \refresh_counter[10] (
	.clk(clk_clk),
	.d(\refresh_counter~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[10]~q ),
	.prn(vcc));
defparam \refresh_counter[10] .is_wysiwyg = "true";
defparam \refresh_counter[10] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~2 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~17_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~2 .extended_lut = "off";
defparam \refresh_counter~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \refresh_counter~2 .shared_arith = "off";

dffeas \refresh_counter[11] (
	.clk(clk_clk),
	.d(\refresh_counter~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[11]~q ),
	.prn(vcc));
defparam \refresh_counter[11] .is_wysiwyg = "true";
defparam \refresh_counter[11] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_counter[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000000000FF00;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \refresh_counter~1 (
	.dataa(!\Equal0~2_combout ),
	.datab(!\Add0~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_counter~1 .extended_lut = "off";
defparam \refresh_counter~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \refresh_counter~1 .shared_arith = "off";

dffeas \refresh_counter[12] (
	.clk(clk_clk),
	.d(\refresh_counter~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[12]~q ),
	.prn(vcc));
defparam \refresh_counter[12] .is_wysiwyg = "true";
defparam \refresh_counter[12] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\refresh_counter[12]~q ),
	.datab(!\refresh_counter[11]~q ),
	.datac(!\refresh_counter[10]~q ),
	.datad(!\refresh_counter[9]~q ),
	.datae(!\refresh_counter[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\refresh_counter[6]~q ),
	.datab(!\refresh_counter[5]~q ),
	.datac(!\refresh_counter[4]~q ),
	.datad(!\refresh_counter[3]~q ),
	.datae(!\refresh_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\refresh_counter[7]~q ),
	.datab(!\refresh_counter[1]~q ),
	.datac(!\refresh_counter[0]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \i_count[1]~0 (
	.dataa(!\i_state.101~q ),
	.datab(!\i_state.000~q ),
	.datac(!\i_state.011~q ),
	.datad(!\i_count[2]~q ),
	.datae(!\i_count[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_count[1]~0 .extended_lut = "off";
defparam \i_count[1]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \i_count[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \i_count[0]~2 (
	.dataa(!\i_state.011~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_count[0]~q ),
	.datad(!\i_count[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_count[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_count[0]~2 .extended_lut = "off";
defparam \i_count[0]~2 .lut_mask = 64'hB77BB77BB77BB77B;
defparam \i_count[0]~2 .shared_arith = "off";

dffeas \i_count[0] (
	.clk(clk_clk),
	.d(\i_count[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[0]~q ),
	.prn(vcc));
defparam \i_count[0] .is_wysiwyg = "true";
defparam \i_count[0] .power_up = "low";

cyclonev_lcell_comb \i_count[1]~1 (
	.dataa(!\i_state.011~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_count[1]~q ),
	.datad(!\i_count[0]~q ),
	.datae(!\i_count[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_count[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_count[1]~1 .extended_lut = "off";
defparam \i_count[1]~1 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \i_count[1]~1 .shared_arith = "off";

dffeas \i_count[1] (
	.clk(clk_clk),
	.d(\i_count[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[1]~q ),
	.prn(vcc));
defparam \i_count[1] .is_wysiwyg = "true";
defparam \i_count[1] .power_up = "low";

cyclonev_lcell_comb WideOr6(
	.dataa(!\i_state.101~q ),
	.datab(!\i_state.000~q ),
	.datac(!\i_state.011~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr6~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr6.extended_lut = "off";
defparam WideOr6.lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam WideOr6.shared_arith = "off";

cyclonev_lcell_comb \i_next.000~0 (
	.dataa(!\i_next.000~q ),
	.datab(!\WideOr6~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_next.000~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_next.000~0 .extended_lut = "off";
defparam \i_next.000~0 .lut_mask = 64'h7777777777777777;
defparam \i_next.000~0 .shared_arith = "off";

dffeas \i_next.000 (
	.clk(clk_clk),
	.d(\i_next.000~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.000~q ),
	.prn(vcc));
defparam \i_next.000 .is_wysiwyg = "true";
defparam \i_next.000 .power_up = "low";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!\i_state.000~q ),
	.datab(!\i_state.011~q ),
	.datac(!\Equal0~2_combout ),
	.datad(!\i_count[2]~q ),
	.datae(!\i_count[1]~q ),
	.dataf(!\i_next.000~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \Selector7~0 .shared_arith = "off";

dffeas \i_state.000 (
	.clk(clk_clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.000~q ),
	.prn(vcc));
defparam \i_state.000 .is_wysiwyg = "true";
defparam \i_state.000 .power_up = "low";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!\i_state.011~q ),
	.datab(!\i_count[1]~q ),
	.datac(!\i_count[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector13~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~1 (
	.dataa(!\i_state.111~q ),
	.datab(!\i_state.101~q ),
	.datac(!\i_state.000~q ),
	.datad(!\i_count[2]~q ),
	.datae(!\Selector13~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~1 .extended_lut = "off";
defparam \Selector13~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \Selector13~1 .shared_arith = "off";

dffeas \i_count[2] (
	.clk(clk_clk),
	.d(\Selector13~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[2]~q ),
	.prn(vcc));
defparam \i_count[2] .is_wysiwyg = "true";
defparam \i_count[2] .power_up = "low";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\i_state.000~q ),
	.datab(!\Equal0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Selector8~0 .shared_arith = "off";

dffeas \i_state.001 (
	.clk(clk_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.001~q ),
	.prn(vcc));
defparam \i_state.001 .is_wysiwyg = "true";
defparam \i_state.001 .power_up = "low";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!\i_state.000~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_refs[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \Selector6~0 .shared_arith = "off";

dffeas \i_refs[0] (
	.clk(clk_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[0]~q ),
	.prn(vcc));
defparam \i_refs[0] .is_wysiwyg = "true";
defparam \i_refs[0] .power_up = "low";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\i_state.000~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_refs[1]~q ),
	.datad(!\i_refs[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \Selector5~0 .shared_arith = "off";

dffeas \i_refs[1] (
	.clk(clk_clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[1]~q ),
	.prn(vcc));
defparam \i_refs[1] .is_wysiwyg = "true";
defparam \i_refs[1] .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!\i_state.000~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_refs[2]~q ),
	.datad(!\i_refs[1]~q ),
	.datae(!\i_refs[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \Selector4~0 .shared_arith = "off";

dffeas \i_refs[2] (
	.clk(clk_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[2]~q ),
	.prn(vcc));
defparam \i_refs[2] .is_wysiwyg = "true";
defparam \i_refs[2] .power_up = "low";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!\i_refs[2]~q ),
	.datab(!\i_refs[1]~q ),
	.datac(!\i_refs[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Selector18~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!\i_state.001~q ),
	.datab(!\i_state.010~q ),
	.datac(!\i_next.010~q ),
	.datad(!\WideOr6~combout ),
	.datae(!\Selector18~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \Selector16~0 .shared_arith = "off";

dffeas \i_next.010 (
	.clk(clk_clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.010~q ),
	.prn(vcc));
defparam \i_next.010 .is_wysiwyg = "true";
defparam \i_next.010 .power_up = "low";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!\i_state.011~q ),
	.datab(!\i_count[2]~q ),
	.datac(!\i_count[1]~q ),
	.datad(!\i_next.010~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \Selector9~0 .shared_arith = "off";

dffeas \i_state.010 (
	.clk(clk_clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.010~q ),
	.prn(vcc));
defparam \i_state.010 .is_wysiwyg = "true";
defparam \i_state.010 .power_up = "low";

cyclonev_lcell_comb \Selector18~1 (
	.dataa(!\i_state.010~q ),
	.datab(!\i_next.111~q ),
	.datac(!\WideOr6~combout ),
	.datad(!\Selector18~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~1 .extended_lut = "off";
defparam \Selector18~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \Selector18~1 .shared_arith = "off";

dffeas \i_next.111 (
	.clk(clk_clk),
	.d(\Selector18~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.111~q ),
	.prn(vcc));
defparam \i_next.111 .is_wysiwyg = "true";
defparam \i_next.111 .power_up = "low";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!\i_state.011~q ),
	.datab(!\i_next.111~q ),
	.datac(!\i_count[2]~q ),
	.datad(!\i_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Selector12~0 .shared_arith = "off";

dffeas \i_state.111 (
	.clk(clk_clk),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.111~q ),
	.prn(vcc));
defparam \i_state.111 .is_wysiwyg = "true";
defparam \i_state.111 .power_up = "low";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!\i_state.111~q ),
	.datab(!\i_state.001~q ),
	.datac(!\i_state.011~q ),
	.datad(!\i_state.010~q ),
	.datae(!\i_count[2]~q ),
	.dataf(!\i_count[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Selector10~0 .shared_arith = "off";

dffeas \i_state.011 (
	.clk(clk_clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.011~q ),
	.prn(vcc));
defparam \i_state.011 .is_wysiwyg = "true";
defparam \i_state.011 .power_up = "low";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\i_state.111~q ),
	.datab(!\i_next.101~q ),
	.datac(!\WideOr6~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Selector17~0 .shared_arith = "off";

dffeas \i_next.101 (
	.clk(clk_clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.101~q ),
	.prn(vcc));
defparam \i_next.101 .is_wysiwyg = "true";
defparam \i_next.101 .power_up = "low";

cyclonev_lcell_comb \i_state.101~0 (
	.dataa(!\i_state.101~q ),
	.datab(!\i_state.011~q ),
	.datac(!\i_count[2]~q ),
	.datad(!\i_count[1]~q ),
	.datae(!\i_next.101~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_state.101~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_state.101~0 .extended_lut = "off";
defparam \i_state.101~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \i_state.101~0 .shared_arith = "off";

dffeas \i_state.101 (
	.clk(clk_clk),
	.d(\i_state.101~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.101~q ),
	.prn(vcc));
defparam \i_state.101 .is_wysiwyg = "true";
defparam \i_state.101 .power_up = "low";

cyclonev_lcell_comb \init_done~0 (
	.dataa(!\init_done~q ),
	.datab(!\i_state.101~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\init_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \init_done~0 .extended_lut = "off";
defparam \init_done~0 .lut_mask = 64'h7777777777777777;
defparam \init_done~0 .shared_arith = "off";

dffeas init_done(
	.clk(clk_clk),
	.d(\init_done~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\init_done~q ),
	.prn(vcc));
defparam init_done.is_wysiwyg = "true";
defparam init_done.power_up = "low";

cyclonev_lcell_comb \Selector32~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\Selector41~0_combout ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_state.100000000~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \Selector32~0 .shared_arith = "off";

dffeas \m_state.100000000 (
	.clk(clk_clk),
	.d(\Selector32~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.100000000~q ),
	.prn(vcc));
defparam \m_state.100000000 .is_wysiwyg = "true";
defparam \m_state.100000000 .power_up = "low";

dffeas \active_addr[14] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[50]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[14]~q ),
	.prn(vcc));
defparam \active_addr[14] .is_wysiwyg = "true";
defparam \active_addr[14] .power_up = "low";

cyclonev_lcell_comb \Equal3~5 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[14]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[50]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[50]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~5 .extended_lut = "off";
defparam \Equal3~5 .lut_mask = 64'h6996699669966996;
defparam \Equal3~5 .shared_arith = "off";

dffeas \active_addr[15] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[51]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[15]~q ),
	.prn(vcc));
defparam \active_addr[15] .is_wysiwyg = "true";
defparam \active_addr[15] .power_up = "low";

cyclonev_lcell_comb \Equal3~6 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[15]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[51]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[51]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~6 .extended_lut = "off";
defparam \Equal3~6 .lut_mask = 64'h6996699669966996;
defparam \Equal3~6 .shared_arith = "off";

dffeas \active_addr[16] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[52]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[16]~q ),
	.prn(vcc));
defparam \active_addr[16] .is_wysiwyg = "true";
defparam \active_addr[16] .power_up = "low";

cyclonev_lcell_comb \Equal3~7 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[16]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[52]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[52]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~7 .extended_lut = "off";
defparam \Equal3~7 .lut_mask = 64'h6996699669966996;
defparam \Equal3~7 .shared_arith = "off";

dffeas \active_addr[17] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[53]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[17]~q ),
	.prn(vcc));
defparam \active_addr[17] .is_wysiwyg = "true";
defparam \active_addr[17] .power_up = "low";

cyclonev_lcell_comb \Equal3~8 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[17]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[53]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[53]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~8 .extended_lut = "off";
defparam \Equal3~8 .lut_mask = 64'h6996699669966996;
defparam \Equal3~8 .shared_arith = "off";

dffeas \active_addr[18] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[54]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[18]~q ),
	.prn(vcc));
defparam \active_addr[18] .is_wysiwyg = "true";
defparam \active_addr[18] .power_up = "low";

cyclonev_lcell_comb \Equal3~9 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[18]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[54]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[54]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~9 .extended_lut = "off";
defparam \Equal3~9 .lut_mask = 64'h6996699669966996;
defparam \Equal3~9 .shared_arith = "off";

dffeas \active_addr[19] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[55]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[19]~q ),
	.prn(vcc));
defparam \active_addr[19] .is_wysiwyg = "true";
defparam \active_addr[19] .power_up = "low";

cyclonev_lcell_comb \Equal3~10 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datab(!\active_addr[19]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[55]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[55]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~10 .extended_lut = "off";
defparam \Equal3~10 .lut_mask = 64'h6996699669966996;
defparam \Equal3~10 .shared_arith = "off";

cyclonev_lcell_comb \pending~3 (
	.dataa(!\Equal3~5_combout ),
	.datab(!\Equal3~6_combout ),
	.datac(!\Equal3~7_combout ),
	.datad(!\Equal3~8_combout ),
	.datae(!\Equal3~9_combout ),
	.dataf(!\Equal3~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending~3 .extended_lut = "off";
defparam \pending~3 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \pending~3 .shared_arith = "off";

cyclonev_lcell_comb \pending~4 (
	.dataa(!\pending~0_combout ),
	.datab(!\pending~2_combout ),
	.datac(!\pending~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending~4 .extended_lut = "off";
defparam \pending~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \pending~4 .shared_arith = "off";

cyclonev_lcell_comb \m_next~17 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_next~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_next~17 .extended_lut = "off";
defparam \m_next~17 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \m_next~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~0 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.100000000~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~0 .extended_lut = "off";
defparam \Selector35~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \Selector35~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~1 (
	.dataa(!\m_state.010000000~q ),
	.datab(!\init_done~q ),
	.datac(!\m_state.000000001~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~1 .extended_lut = "off";
defparam \Selector35~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Selector35~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector34~0 (
	.dataa(!\active_rnw~q ),
	.datab(!\m_state.000000010~q ),
	.datac(!\m_next.000001000~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~0 .extended_lut = "off";
defparam \Selector34~0 .lut_mask = 64'h4747474747474747;
defparam \Selector34~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector34~1 (
	.dataa(!\m_state.100000000~q ),
	.datab(!\m_next~17_combout ),
	.datac(!\Selector35~0_combout ),
	.datad(!\Selector35~1_combout ),
	.datae(!\Selector34~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~1 .extended_lut = "off";
defparam \Selector34~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Selector34~1 .shared_arith = "off";

dffeas \m_next.000001000 (
	.clk(clk_clk),
	.d(\Selector34~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000001000~q ),
	.prn(vcc));
defparam \m_next.000001000 .is_wysiwyg = "true";
defparam \m_next.000001000 .power_up = "low";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\m_state.100000000~q ),
	.datac(!\refresh_request~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~1 (
	.dataa(!\pending~0_combout ),
	.datab(!\pending~2_combout ),
	.datac(!\pending~3_combout ),
	.datad(!\refresh_request~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~1 .extended_lut = "off";
defparam \Selector28~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Selector28~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!\m_state.100000000~q ),
	.datab(!\m_state.000100000~q ),
	.datac(!\refresh_request~q ),
	.datad(!\m_count[1]~q ),
	.datae(!\m_next~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \Selector29~0 .shared_arith = "off";

dffeas \m_state.000100000 (
	.clk(clk_clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000100000~q ),
	.prn(vcc));
defparam \m_state.000100000 .is_wysiwyg = "true";
defparam \m_state.000100000 .power_up = "low";

cyclonev_lcell_comb \Selector24~1 (
	.dataa(!\m_state.000100000~q ),
	.datab(!\m_count[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~1 .extended_lut = "off";
defparam \Selector24~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector24~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector30~1 (
	.dataa(!\Selector30~0_combout ),
	.datab(!\refresh_request~q ),
	.datac(!\Selector24~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector30~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector30~1 .extended_lut = "off";
defparam \Selector30~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector30~1 .shared_arith = "off";

dffeas \m_state.001000000 (
	.clk(clk_clk),
	.d(\Selector30~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.001000000~q ),
	.prn(vcc));
defparam \m_state.001000000 .is_wysiwyg = "true";
defparam \m_state.001000000 .power_up = "low";

cyclonev_lcell_comb \Selector36~2 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~4_combout ),
	.datac(!\m_state.001000000~q ),
	.datad(!\m_state.100000000~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~2 .extended_lut = "off";
defparam \Selector36~2 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Selector36~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~3 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~0_combout ),
	.datac(!\pending~2_combout ),
	.datad(!\pending~3_combout ),
	.datae(!\WideOr9~0_combout ),
	.dataf(!\WideOr8~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~3 .extended_lut = "off";
defparam \Selector28~3 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \Selector28~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~4 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\init_done~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~4 .extended_lut = "off";
defparam \Selector28~4 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \Selector28~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~5 (
	.dataa(!\Selector24~1_combout ),
	.datab(!\Selector28~3_combout ),
	.datac(!\Selector28~4_combout ),
	.datad(!\Selector28~0_combout ),
	.datae(!\Selector28~1_combout ),
	.dataf(!\Selector24~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~5 .extended_lut = "off";
defparam \Selector28~5 .lut_mask = 64'hFFFFFFFF6996FFFF;
defparam \Selector28~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~2 (
	.dataa(!\active_rnw~q ),
	.datab(!\m_state.000000010~q ),
	.datac(!\m_next.000010000~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~2 .extended_lut = "off";
defparam \Selector35~2 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \Selector35~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~3 (
	.dataa(!\m_state.100000000~q ),
	.datab(!\m_next~17_combout ),
	.datac(!\Selector35~0_combout ),
	.datad(!\Selector35~1_combout ),
	.datae(!\Selector35~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~3 .extended_lut = "off";
defparam \Selector35~3 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Selector35~3 .shared_arith = "off";

dffeas \m_next.000010000 (
	.clk(clk_clk),
	.d(\Selector35~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000010000~q ),
	.prn(vcc));
defparam \m_next.000010000 .is_wysiwyg = "true";
defparam \m_next.000010000 .power_up = "low";

cyclonev_lcell_comb \Selector28~6 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_data[61]~19_combout ),
	.datab(!\m_state.000010000~q ),
	.datac(!\Selector28~2_combout ),
	.datad(!\Selector28~5_combout ),
	.datae(!\m_next.000010000~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~6 .extended_lut = "off";
defparam \Selector28~6 .lut_mask = 64'hBFFBFFFFBFFBFFFF;
defparam \Selector28~6 .shared_arith = "off";

dffeas \m_state.000010000 (
	.clk(clk_clk),
	.d(\Selector28~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000010000~q ),
	.prn(vcc));
defparam \m_state.000010000 .is_wysiwyg = "true";
defparam \m_state.000010000 .power_up = "low";

cyclonev_lcell_comb \Selector38~0 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\m_state.000010000~q ),
	.datac(!\refresh_request~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~0 .extended_lut = "off";
defparam \Selector38~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Selector38~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector38~1 (
	.dataa(!\m_state.000001000~q ),
	.datab(!\init_done~q ),
	.datac(!\m_state.000000001~q ),
	.datad(!\refresh_request~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~1 .extended_lut = "off";
defparam \Selector38~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Selector38~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~4_combout ),
	.datac(!\m_state.000010000~q ),
	.datad(!\m_state.100000000~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~0 .extended_lut = "off";
defparam \Selector39~0 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \Selector39~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~1 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\m_state.000001000~q ),
	.datac(!\Selector30~0_combout ),
	.datad(!\refresh_request~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~1 .extended_lut = "off";
defparam \Selector39~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector39~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~2 (
	.dataa(!\m_state.000000100~q ),
	.datab(!\m_state.000100000~q ),
	.datac(!\m_count[1]~q ),
	.datad(!\m_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~2 .extended_lut = "off";
defparam \Selector39~2 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \Selector39~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~3 (
	.dataa(!\m_state.000001000~q ),
	.datab(!\m_state.001000000~q ),
	.datac(!\m_state.000000001~q ),
	.datad(!\Selector39~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~3 .extended_lut = "off";
defparam \Selector39~3 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \Selector39~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~4 (
	.dataa(!\m_state.000000100~q ),
	.datab(!\m_state.000100000~q ),
	.datac(!\m_count[1]~q ),
	.datad(!\m_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~4 .extended_lut = "off";
defparam \Selector39~4 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \Selector39~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector39~5 (
	.dataa(!\Selector39~0_combout ),
	.datab(!\Selector39~1_combout ),
	.datac(!\Selector39~3_combout ),
	.datad(!\Selector39~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~5 .extended_lut = "off";
defparam \Selector39~5 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Selector39~5 .shared_arith = "off";

dffeas \m_count[0] (
	.clk(clk_clk),
	.d(\Selector39~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[0]~q ),
	.prn(vcc));
defparam \m_count[0] .is_wysiwyg = "true";
defparam \m_count[0] .power_up = "low";

cyclonev_lcell_comb \Selector38~2 (
	.dataa(!\m_state.000000100~q ),
	.datab(!\m_state.000100000~q ),
	.datac(!\m_count[1]~q ),
	.datad(!\m_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~2 .extended_lut = "off";
defparam \Selector38~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector38~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector38~3 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\m_state.000001000~q ),
	.datac(!\m_state.010000000~q ),
	.datad(!\refresh_request~q ),
	.datae(!\Selector38~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~3 .extended_lut = "off";
defparam \Selector38~3 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Selector38~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector38~4 (
	.dataa(!\m_count[1]~q ),
	.datab(!\Selector36~2_combout ),
	.datac(!\Selector38~0_combout ),
	.datad(!\Selector38~1_combout ),
	.datae(!\Selector38~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~4 .extended_lut = "off";
defparam \Selector38~4 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \Selector38~4 .shared_arith = "off";

dffeas \m_count[1] (
	.clk(clk_clk),
	.d(\Selector38~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[1]~q ),
	.prn(vcc));
defparam \m_count[1] .is_wysiwyg = "true";
defparam \m_count[1] .power_up = "low";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!\m_state.000000100~q ),
	.datab(!\m_count[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~2 (
	.dataa(!\Selector28~0_combout ),
	.datab(!\Selector28~1_combout ),
	.datac(!\Selector24~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~2 .extended_lut = "off";
defparam \Selector28~2 .lut_mask = 64'hD8D8D8D8D8D8D8D8;
defparam \Selector28~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|rd_data[61]~19_combout ),
	.datab(!\m_state.000001000~q ),
	.datac(!\m_next.000001000~q ),
	.datad(!\Selector28~2_combout ),
	.datae(!\Selector28~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \Selector27~0 .shared_arith = "off";

dffeas \m_state.000001000 (
	.clk(clk_clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000001000~q ),
	.prn(vcc));
defparam \m_state.000001000 .is_wysiwyg = "true";
defparam \m_state.000001000 .power_up = "low";

cyclonev_lcell_comb \WideOr9~0 (
	.dataa(!\m_state.000001000~q ),
	.datab(!\m_state.000010000~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr9~0 .extended_lut = "off";
defparam \WideOr9~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \WideOr9~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!\m_state.100000000~q ),
	.datab(!\m_state.000000100~q ),
	.datac(!\refresh_request~q ),
	.datad(!\WideOr8~0_combout ),
	.datae(!\m_count[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.000000100~q ),
	.datad(!\refresh_request~q ),
	.datae(!\Selector26~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \Selector26~1 .shared_arith = "off";

dffeas \m_state.000000100 (
	.clk(clk_clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000100~q ),
	.prn(vcc));
defparam \m_state.000000100 .is_wysiwyg = "true";
defparam \m_state.000000100 .power_up = "low";

cyclonev_lcell_comb \Selector36~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~4_combout ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_state.001000000~q ),
	.datae(!\m_state.100000000~q ),
	.dataf(!\refresh_request~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~0 .extended_lut = "off";
defparam \Selector36~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \Selector36~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector36~1 (
	.dataa(!\Selector30~0_combout ),
	.datab(!\m_state.000000100~q ),
	.datac(!\m_state.000100000~q ),
	.datad(!\refresh_request~q ),
	.datae(!\m_next.010000000~q ),
	.dataf(!\Selector36~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~1 .extended_lut = "off";
defparam \Selector36~1 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \Selector36~1 .shared_arith = "off";

dffeas \m_next.010000000 (
	.clk(clk_clk),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.010000000~q ),
	.prn(vcc));
defparam \m_next.010000000 .is_wysiwyg = "true";
defparam \m_next.010000000 .power_up = "low";

cyclonev_lcell_comb \Selector24~2 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\m_state.100000000~q ),
	.datac(!\init_done~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~2 .extended_lut = "off";
defparam \Selector24~2 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \Selector24~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~3 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\refresh_request~q ),
	.datad(!\WideOr8~0_combout ),
	.datae(!\Selector24~1_combout ),
	.dataf(!\Selector24~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~3 .extended_lut = "off";
defparam \Selector24~3 .lut_mask = 64'h6996966996696996;
defparam \Selector24~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector31~0 (
	.dataa(!\m_next.010000000~q ),
	.datab(!\Selector24~0_combout ),
	.datac(!\Selector24~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector31~0 .extended_lut = "off";
defparam \Selector31~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector31~0 .shared_arith = "off";

dffeas \m_state.010000000 (
	.clk(clk_clk),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.010000000~q ),
	.prn(vcc));
defparam \m_state.010000000 .is_wysiwyg = "true";
defparam \m_state.010000000 .power_up = "low";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!\m_state.010000000~q ),
	.datab(!\init_done~q ),
	.datac(!\m_state.000000001~q ),
	.datad(!\ack_refresh_request~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Selector23~0 .shared_arith = "off";

dffeas ack_refresh_request(
	.clk(clk_clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ack_refresh_request~q ),
	.prn(vcc));
defparam ack_refresh_request.is_wysiwyg = "true";
defparam ack_refresh_request.power_up = "low";

cyclonev_lcell_comb \refresh_request~0 (
	.dataa(!\init_done~q ),
	.datab(!\refresh_request~q ),
	.datac(!\ack_refresh_request~q ),
	.datad(!\Equal0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_request~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_request~0 .extended_lut = "off";
defparam \refresh_request~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \refresh_request~0 .shared_arith = "off";

dffeas refresh_request(
	.clk(clk_clk),
	.d(\refresh_request~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_request~q ),
	.prn(vcc));
defparam refresh_request.is_wysiwyg = "true";
defparam refresh_request.power_up = "low";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\Selector30~0_combout ),
	.datac(!\refresh_request~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Selector25~0 .shared_arith = "off";

dffeas \m_state.000000010 (
	.clk(clk_clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000010~q ),
	.prn(vcc));
defparam \m_state.000000010 .is_wysiwyg = "true";
defparam \m_state.000000010 .power_up = "low";

cyclonev_lcell_comb \WideOr8~0 (
	.dataa(!\m_state.000000010~q ),
	.datab(!\m_state.001000000~q ),
	.datac(!\m_state.010000000~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr8~0 .extended_lut = "off";
defparam \WideOr8~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \WideOr8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~0 (
	.dataa(!\m_state.001000000~q ),
	.datab(!\m_state.000000001~q ),
	.datac(!\m_state.000000100~q ),
	.datad(!\m_state.000100000~q ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \Selector33~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~1 (
	.dataa(!\WideOr9~0_combout ),
	.datab(!\m_state.100000000~q ),
	.datac(!\m_next.000000001~q ),
	.datad(!\Selector35~1_combout ),
	.datae(!\Selector33~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~1 .extended_lut = "off";
defparam \Selector33~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \Selector33~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector33~2 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~4_combout ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_state.100000000~q ),
	.datae(!\refresh_request~q ),
	.dataf(!\Selector33~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~2 .extended_lut = "off";
defparam \Selector33~2 .lut_mask = 64'hFF7FDF5FFFFFFFFF;
defparam \Selector33~2 .shared_arith = "off";

dffeas \m_next.000000001 (
	.clk(clk_clk),
	.d(\Selector33~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000000001~q ),
	.prn(vcc));
defparam \m_next.000000001 .is_wysiwyg = "true";
defparam \m_next.000000001 .power_up = "low";

cyclonev_lcell_comb \Selector24~4 (
	.dataa(!\init_done~q ),
	.datab(!\m_state.000000001~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\Selector24~0_combout ),
	.datae(!\Selector24~3_combout ),
	.dataf(!\m_next.000000001~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~4 .extended_lut = "off";
defparam \Selector24~4 .lut_mask = 64'hF7FFFFF7FFFFFFFF;
defparam \Selector24~4 .shared_arith = "off";

dffeas \m_state.000000001 (
	.clk(clk_clk),
	.d(\Selector24~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000001~q ),
	.prn(vcc));
defparam \m_state.000000001 .is_wysiwyg = "true";
defparam \m_state.000000001 .power_up = "low";

cyclonev_lcell_comb \Selector30~0 (
	.dataa(!\init_done~q ),
	.datab(!\m_state.000000001~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector30~0 .extended_lut = "off";
defparam \Selector30~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector30~0 .shared_arith = "off";

cyclonev_lcell_comb \active_cs_n~0 (
	.dataa(!r_sync_rst),
	.datab(!\active_cs_n~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(!\Selector30~0_combout ),
	.datae(!\refresh_request~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\active_cs_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \active_cs_n~0 .extended_lut = "off";
defparam \active_cs_n~0 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \active_cs_n~0 .shared_arith = "off";

dffeas active_cs_n(
	.clk(clk_clk),
	.d(\active_cs_n~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\active_cs_n~q ),
	.prn(vcc));
defparam active_cs_n.is_wysiwyg = "true";
defparam active_cs_n.power_up = "low";

cyclonev_lcell_comb \pending~1 (
	.dataa(!\active_rnw~q ),
	.datab(!\the_sdram_demo_sdram_input_efifo_module|rd_address~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|entry_1[61]~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|entry_0[61]~q ),
	.datae(!\active_cs_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending~1 .extended_lut = "off";
defparam \pending~1 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \pending~1 .shared_arith = "off";

cyclonev_lcell_comb \pending~2 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal2~1_combout ),
	.datac(!\Equal3~2_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(!\Equal3~4_combout ),
	.dataf(!\pending~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending~2 .extended_lut = "off";
defparam \pending~2 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \pending~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector41~0 (
	.dataa(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(!\pending~0_combout ),
	.datac(!\pending~2_combout ),
	.datad(!\pending~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector41~0 .extended_lut = "off";
defparam \Selector41~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Selector41~0 .shared_arith = "off";

cyclonev_lcell_comb \active_rnw~0 (
	.dataa(!entries_1),
	.datab(!entries_0),
	.datac(!\init_done~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\active_rnw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \active_rnw~0 .extended_lut = "off";
defparam \active_rnw~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \active_rnw~0 .shared_arith = "off";

cyclonev_lcell_comb \active_rnw~1 (
	.dataa(!r_sync_rst),
	.datab(!\refresh_request~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\active_rnw~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \active_rnw~1 .extended_lut = "off";
defparam \active_rnw~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \active_rnw~1 .shared_arith = "off";

cyclonev_lcell_comb \active_rnw~2 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.100000000~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\active_rnw~0_combout ),
	.dataf(!\active_rnw~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\active_rnw~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \active_rnw~2 .extended_lut = "off";
defparam \active_rnw~2 .lut_mask = 64'hCF5FFFFFFFFFFFFF;
defparam \active_rnw~2 .shared_arith = "off";

dffeas \active_addr[0] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[36]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[0]~q ),
	.prn(vcc));
defparam \active_addr[0] .is_wysiwyg = "true";
defparam \active_addr[0] .power_up = "low";

cyclonev_lcell_comb \Selector41~1 (
	.dataa(!\Selector41~0_combout ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.100000000~q ),
	.datad(!\refresh_request~q ),
	.datae(!\Selector25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector41~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector41~1 .extended_lut = "off";
defparam \Selector41~1 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \Selector41~1 .shared_arith = "off";

dffeas f_pop(
	.clk(clk_clk),
	.d(\Selector41~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\f_pop~q ),
	.prn(vcc));
defparam f_pop.is_wysiwyg = "true";
defparam f_pop.power_up = "low";

cyclonev_lcell_comb \m_addr[6]~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_state.000000010~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_addr[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_addr[6]~0 .extended_lut = "off";
defparam \m_addr[6]~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \m_addr[6]~0 .shared_arith = "off";

dffeas \i_addr[12] (
	.clk(clk_clk),
	.d(\i_state.111~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_addr[12]~q ),
	.prn(vcc));
defparam \i_addr[12] .is_wysiwyg = "true";
defparam \i_addr[12] .power_up = "low";

cyclonev_lcell_comb \Selector116~0 (
	.dataa(!\active_addr[0]~q ),
	.datab(!\active_addr[11]~q ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_addr[6]~0_combout ),
	.datae(!\the_sdram_demo_sdram_input_efifo_module|rd_data[36]~2_combout ),
	.dataf(!\i_addr[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector116~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector116~0 .extended_lut = "off";
defparam \Selector116~0 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \Selector116~0 .shared_arith = "off";

cyclonev_lcell_comb \m_addr[6]~1 (
	.dataa(!\m_state.010000000~q ),
	.datab(!\m_state.100000000~q ),
	.datac(!\Selector30~0_combout ),
	.datad(!\m_state.000000100~q ),
	.datae(!\m_state.000100000~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_addr[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_addr[6]~1 .extended_lut = "off";
defparam \m_addr[6]~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \m_addr[6]~1 .shared_arith = "off";

dffeas \active_addr[1] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[37]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[1]~q ),
	.prn(vcc));
defparam \active_addr[1] .is_wysiwyg = "true";
defparam \active_addr[1] .power_up = "low";

cyclonev_lcell_comb \Selector115~0 (
	.dataa(!\active_addr[12]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[1]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[37]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector115~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector115~0 .extended_lut = "off";
defparam \Selector115~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector115~0 .shared_arith = "off";

dffeas \active_addr[2] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[38]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[2]~q ),
	.prn(vcc));
defparam \active_addr[2] .is_wysiwyg = "true";
defparam \active_addr[2] .power_up = "low";

cyclonev_lcell_comb \Selector114~0 (
	.dataa(!\active_addr[13]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[2]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[38]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector114~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector114~0 .extended_lut = "off";
defparam \Selector114~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector114~0 .shared_arith = "off";

dffeas \active_addr[3] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[39]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[3]~q ),
	.prn(vcc));
defparam \active_addr[3] .is_wysiwyg = "true";
defparam \active_addr[3] .power_up = "low";

cyclonev_lcell_comb \Selector113~0 (
	.dataa(!\active_addr[14]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[3]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[39]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector113~0 .extended_lut = "off";
defparam \Selector113~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector113~0 .shared_arith = "off";

dffeas \active_addr[6] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[42]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[6]~q ),
	.prn(vcc));
defparam \active_addr[6] .is_wysiwyg = "true";
defparam \active_addr[6] .power_up = "low";

cyclonev_lcell_comb \Selector110~0 (
	.dataa(!\active_addr[17]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[6]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[42]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector110~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector110~0 .extended_lut = "off";
defparam \Selector110~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector110~0 .shared_arith = "off";

dffeas \active_addr[7] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[43]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[7]~q ),
	.prn(vcc));
defparam \active_addr[7] .is_wysiwyg = "true";
defparam \active_addr[7] .power_up = "low";

cyclonev_lcell_comb \Selector109~0 (
	.dataa(!\active_addr[18]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[7]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[43]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector109~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector109~0 .extended_lut = "off";
defparam \Selector109~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector109~0 .shared_arith = "off";

dffeas \active_addr[8] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[44]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[8]~q ),
	.prn(vcc));
defparam \active_addr[8] .is_wysiwyg = "true";
defparam \active_addr[8] .power_up = "low";

cyclonev_lcell_comb \Selector108~0 (
	.dataa(!\active_addr[19]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[8]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[44]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector108~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector108~0 .extended_lut = "off";
defparam \Selector108~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector108~0 .shared_arith = "off";

dffeas \active_addr[9] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[45]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[9]~q ),
	.prn(vcc));
defparam \active_addr[9] .is_wysiwyg = "true";
defparam \active_addr[9] .power_up = "low";

cyclonev_lcell_comb \Selector107~0 (
	.dataa(!\active_addr[20]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_addr[6]~0_combout ),
	.datad(!\i_addr[12]~q ),
	.datae(!\active_addr[9]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[45]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector107~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector107~0 .extended_lut = "off";
defparam \Selector107~0 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \Selector107~0 .shared_arith = "off";

cyclonev_lcell_comb \always5~0 (
	.dataa(!\f_pop~q ),
	.datab(!\the_sdram_demo_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(!\pending~0_combout ),
	.datad(!\pending~2_combout ),
	.datae(!\pending~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \always5~0 .shared_arith = "off";

dffeas \active_addr[4] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[40]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[4]~q ),
	.prn(vcc));
defparam \active_addr[4] .is_wysiwyg = "true";
defparam \active_addr[4] .power_up = "low";

cyclonev_lcell_comb \Selector112~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\WideOr9~0_combout ),
	.datad(!\m_state.000000010~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector112~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector112~0 .extended_lut = "off";
defparam \Selector112~0 .lut_mask = 64'hF737F737F737F737;
defparam \Selector112~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector112~1 (
	.dataa(!\active_addr[15]~q ),
	.datab(!\m_addr[6]~0_combout ),
	.datac(!\m_state.001000000~q ),
	.datad(!\active_addr[4]~q ),
	.datae(!\Selector112~0_combout ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[40]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector112~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector112~1 .extended_lut = "off";
defparam \Selector112~1 .lut_mask = 64'h7FFFDFFFFFFFFFFF;
defparam \Selector112~1 .shared_arith = "off";

dffeas \active_addr[5] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[41]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[5]~q ),
	.prn(vcc));
defparam \active_addr[5] .is_wysiwyg = "true";
defparam \active_addr[5] .power_up = "low";

cyclonev_lcell_comb \Selector111~0 (
	.dataa(!\active_addr[16]~q ),
	.datab(!\m_addr[6]~0_combout ),
	.datac(!\m_state.001000000~q ),
	.datad(!\Selector112~0_combout ),
	.datae(!\active_addr[5]~q ),
	.dataf(!\the_sdram_demo_sdram_input_efifo_module|rd_data[41]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector111~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector111~0 .extended_lut = "off";
defparam \Selector111~0 .lut_mask = 64'h7FDFFFFFFFFFFFFF;
defparam \Selector111~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector106~0 (
	.dataa(!\active_addr[21]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\i_addr[12]~q ),
	.datae(!\m_state.001000000~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector106~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector106~0 .extended_lut = "off";
defparam \Selector106~0 .lut_mask = 64'hF737FFFFF737FFFF;
defparam \Selector106~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector105~0 (
	.dataa(!\active_addr[22]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\i_addr[12]~q ),
	.datae(!\m_state.001000000~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector105~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector105~0 .extended_lut = "off";
defparam \Selector105~0 .lut_mask = 64'hF737FFFFF737FFFF;
defparam \Selector105~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector104~0 (
	.dataa(!\active_addr[23]~q ),
	.datab(!\WideOr9~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\i_addr[12]~q ),
	.datae(!\m_state.001000000~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector104~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector104~0 .extended_lut = "off";
defparam \Selector104~0 .lut_mask = 64'hF737FFFFF737FFFF;
defparam \Selector104~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector118~0 (
	.dataa(!\f_pop~q ),
	.datab(!\active_addr[10]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|rd_data[46]~12_combout ),
	.datad(!\Selector41~0_combout ),
	.datae(!\m_state.000000010~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector118~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector118~0 .extended_lut = "off";
defparam \Selector118~0 .lut_mask = 64'hBF7F7FBFBF7F7FBF;
defparam \Selector118~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr16~0 (
	.dataa(!\WideOr9~0_combout ),
	.datab(!\m_state.000000010~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr16~0 .extended_lut = "off";
defparam \WideOr16~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \WideOr16~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector117~0 (
	.dataa(!\f_pop~q ),
	.datab(!\active_addr[24]~q ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|rd_data[60]~13_combout ),
	.datad(!\Selector41~0_combout ),
	.datae(!\m_state.000000010~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector117~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector117~0 .extended_lut = "off";
defparam \Selector117~0 .lut_mask = 64'hBF7F7FBFBF7F7FBF;
defparam \Selector117~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\i_cmd[1]~q ),
	.datab(!\i_state.101~q ),
	.datac(!\i_state.001~q ),
	.datad(!\i_state.000~q ),
	.datae(!\i_state.011~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \Selector2~0 .shared_arith = "off";

dffeas \i_cmd[1] (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[1]~q ),
	.prn(vcc));
defparam \i_cmd[1] .is_wysiwyg = "true";
defparam \i_cmd[1] .power_up = "low";

cyclonev_lcell_comb \Selector21~0 (
	.dataa(!\WideOr9~0_combout ),
	.datab(!\m_state.010000000~q ),
	.datac(!\init_done~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\always5~0_combout ),
	.dataf(!\i_cmd[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \Selector21~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\i_cmd[3]~q ),
	.datab(!\i_state.101~q ),
	.datac(!\i_state.000~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \i_cmd[3] (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[3]~q ),
	.prn(vcc));
defparam \i_cmd[3] .is_wysiwyg = "true";
defparam \i_cmd[3] .power_up = "low";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!\m_state.001000000~q ),
	.datab(!\m_state.010000000~q ),
	.datac(!\m_state.000000001~q ),
	.datad(!\m_state.000000100~q ),
	.datae(!\refresh_request~q ),
	.dataf(!\m_next.010000000~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'hFFFFFFFFFFFFDFEF;
defparam \Selector19~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~1 (
	.dataa(!\active_cs_n~q ),
	.datab(!\init_done~q ),
	.datac(!\m_state.000000001~q ),
	.datad(!\i_cmd[3]~q ),
	.datae(!\refresh_request~q ),
	.dataf(!\Selector19~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~1 .extended_lut = "off";
defparam \Selector19~1 .lut_mask = 64'hBFFFFFFF8FFFFFFF;
defparam \Selector19~1 .shared_arith = "off";

dffeas \active_dqm[0] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[32]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[0]~q ),
	.prn(vcc));
defparam \active_dqm[0] .is_wysiwyg = "true";
defparam \active_dqm[0] .power_up = "low";

cyclonev_lcell_comb \Selector154~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[32]~14_combout ),
	.datae(!\active_dqm[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector154~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector154~0 .extended_lut = "off";
defparam \Selector154~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector154~0 .shared_arith = "off";

dffeas \active_dqm[1] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[33]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[1]~q ),
	.prn(vcc));
defparam \active_dqm[1] .is_wysiwyg = "true";
defparam \active_dqm[1] .power_up = "low";

cyclonev_lcell_comb \Selector153~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[33]~15_combout ),
	.datae(!\active_dqm[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~0 .extended_lut = "off";
defparam \Selector153~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector153~0 .shared_arith = "off";

dffeas \active_dqm[2] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[34]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[2]~q ),
	.prn(vcc));
defparam \active_dqm[2] .is_wysiwyg = "true";
defparam \active_dqm[2] .power_up = "low";

cyclonev_lcell_comb \Selector152~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[34]~16_combout ),
	.datae(!\active_dqm[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~0 .extended_lut = "off";
defparam \Selector152~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector152~0 .shared_arith = "off";

dffeas \active_dqm[3] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[35]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[3]~q ),
	.prn(vcc));
defparam \active_dqm[3] .is_wysiwyg = "true";
defparam \active_dqm[3] .power_up = "low";

cyclonev_lcell_comb \Selector151~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\m_state.000000010~q ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[35]~17_combout ),
	.datae(!\active_dqm[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector151~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector151~0 .extended_lut = "off";
defparam \Selector151~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector151~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\i_cmd[2]~q ),
	.datab(!\i_state.101~q ),
	.datac(!\i_state.000~q ),
	.datad(!\i_state.011~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \Selector1~0 .shared_arith = "off";

dffeas \i_cmd[2] (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[2]~q ),
	.prn(vcc));
defparam \i_cmd[2] .is_wysiwyg = "true";
defparam \i_cmd[2] .power_up = "low";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!\init_done~q ),
	.datab(!\m_state.000000001~q ),
	.datac(!\WideOr8~0_combout ),
	.datad(!\i_cmd[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'hB8FFB8FFB8FFB8FF;
defparam \Selector20~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\i_cmd[0]~q ),
	.datab(!\i_state.101~q ),
	.datac(!\i_state.000~q ),
	.datad(!\i_state.011~q ),
	.datae(!\i_state.010~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \Selector3~0 .shared_arith = "off";

dffeas \i_cmd[0] (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[0]~q ),
	.prn(vcc));
defparam \i_cmd[0] .is_wysiwyg = "true";
defparam \i_cmd[0] .power_up = "low";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!\m_state.000010000~q ),
	.datab(!\m_state.001000000~q ),
	.datac(!\init_done~q ),
	.datad(!\m_state.000000001~q ),
	.datae(!\always5~0_combout ),
	.dataf(!\i_cmd[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'hF7FBFFFFFFFFFFFF;
defparam \Selector22~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!m_cmd_1),
	.datab(!m_cmd_2),
	.datac(!m_cmd_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Equal4~0 .shared_arith = "off";

dffeas \rd_valid[0] (
	.clk(clk_clk),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[0]~q ),
	.prn(vcc));
defparam \rd_valid[0] .is_wysiwyg = "true";
defparam \rd_valid[0] .power_up = "low";

dffeas \rd_valid[1] (
	.clk(clk_clk),
	.d(\rd_valid[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[1]~q ),
	.prn(vcc));
defparam \rd_valid[1] .is_wysiwyg = "true";
defparam \rd_valid[1] .power_up = "low";

dffeas \rd_valid[2] (
	.clk(clk_clk),
	.d(\rd_valid[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[2]~q ),
	.prn(vcc));
defparam \rd_valid[2] .is_wysiwyg = "true";
defparam \rd_valid[2] .power_up = "low";

cyclonev_lcell_comb \m_data[1]~0 (
	.dataa(!\f_pop~q ),
	.datab(!\Selector41~0_combout ),
	.datac(!\m_state.000010000~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_data[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_data[1]~0 .extended_lut = "off";
defparam \m_data[1]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \m_data[1]~0 .shared_arith = "off";

dffeas \active_data[0] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[0]~q ),
	.prn(vcc));
defparam \active_data[0] .is_wysiwyg = "true";
defparam \active_data[0] .power_up = "low";

cyclonev_lcell_comb \WideOr17~0 (
	.dataa(!\m_state.000010000~q ),
	.datab(!\m_state.000000010~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~0 .extended_lut = "off";
defparam \WideOr17~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \WideOr17~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector150~0 (
	.dataa(!m_data_0),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\the_sdram_demo_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.datad(!\active_data[0]~q ),
	.datae(!\WideOr17~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector150~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector150~0 .extended_lut = "off";
defparam \Selector150~0 .lut_mask = 64'h7FFFDFFF7FFFDFFF;
defparam \Selector150~0 .shared_arith = "off";

dffeas \active_data[1] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[1]~q ),
	.prn(vcc));
defparam \active_data[1] .is_wysiwyg = "true";
defparam \active_data[1] .power_up = "low";

cyclonev_lcell_comb \Selector149~0 (
	.dataa(!m_data_1),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.datae(!\active_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector149~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector149~0 .extended_lut = "off";
defparam \Selector149~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector149~0 .shared_arith = "off";

dffeas \active_data[2] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[2]~q ),
	.prn(vcc));
defparam \active_data[2] .is_wysiwyg = "true";
defparam \active_data[2] .power_up = "low";

cyclonev_lcell_comb \Selector148~0 (
	.dataa(!m_data_2),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.datae(!\active_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector148~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector148~0 .extended_lut = "off";
defparam \Selector148~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector148~0 .shared_arith = "off";

dffeas \active_data[3] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[3]~q ),
	.prn(vcc));
defparam \active_data[3] .is_wysiwyg = "true";
defparam \active_data[3] .power_up = "low";

cyclonev_lcell_comb \Selector147~0 (
	.dataa(!m_data_3),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.datae(!\active_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector147~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector147~0 .extended_lut = "off";
defparam \Selector147~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector147~0 .shared_arith = "off";

dffeas \active_data[4] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[4]~q ),
	.prn(vcc));
defparam \active_data[4] .is_wysiwyg = "true";
defparam \active_data[4] .power_up = "low";

cyclonev_lcell_comb \Selector146~0 (
	.dataa(!m_data_4),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.datae(!\active_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector146~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector146~0 .extended_lut = "off";
defparam \Selector146~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector146~0 .shared_arith = "off";

dffeas \active_data[5] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[5]~q ),
	.prn(vcc));
defparam \active_data[5] .is_wysiwyg = "true";
defparam \active_data[5] .power_up = "low";

cyclonev_lcell_comb \Selector145~0 (
	.dataa(!m_data_5),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.datae(!\active_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector145~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector145~0 .extended_lut = "off";
defparam \Selector145~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector145~0 .shared_arith = "off";

dffeas \active_data[6] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[6]~q ),
	.prn(vcc));
defparam \active_data[6] .is_wysiwyg = "true";
defparam \active_data[6] .power_up = "low";

cyclonev_lcell_comb \Selector144~0 (
	.dataa(!m_data_6),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.datae(!\active_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector144~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector144~0 .extended_lut = "off";
defparam \Selector144~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector144~0 .shared_arith = "off";

dffeas \active_data[7] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[7]~q ),
	.prn(vcc));
defparam \active_data[7] .is_wysiwyg = "true";
defparam \active_data[7] .power_up = "low";

cyclonev_lcell_comb \Selector143~0 (
	.dataa(!m_data_7),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.datae(!\active_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector143~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector143~0 .extended_lut = "off";
defparam \Selector143~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector143~0 .shared_arith = "off";

dffeas \active_data[8] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[8]~q ),
	.prn(vcc));
defparam \active_data[8] .is_wysiwyg = "true";
defparam \active_data[8] .power_up = "low";

cyclonev_lcell_comb \Selector142~0 (
	.dataa(!m_data_8),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.datae(!\active_data[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector142~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector142~0 .extended_lut = "off";
defparam \Selector142~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector142~0 .shared_arith = "off";

dffeas \active_data[9] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[9]~q ),
	.prn(vcc));
defparam \active_data[9] .is_wysiwyg = "true";
defparam \active_data[9] .power_up = "low";

cyclonev_lcell_comb \Selector141~0 (
	.dataa(!m_data_9),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.datae(!\active_data[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector141~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector141~0 .extended_lut = "off";
defparam \Selector141~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector141~0 .shared_arith = "off";

dffeas \active_data[10] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[10]~q ),
	.prn(vcc));
defparam \active_data[10] .is_wysiwyg = "true";
defparam \active_data[10] .power_up = "low";

cyclonev_lcell_comb \Selector140~0 (
	.dataa(!m_data_10),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.datae(!\active_data[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector140~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector140~0 .extended_lut = "off";
defparam \Selector140~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector140~0 .shared_arith = "off";

dffeas \active_data[11] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[11]~q ),
	.prn(vcc));
defparam \active_data[11] .is_wysiwyg = "true";
defparam \active_data[11] .power_up = "low";

cyclonev_lcell_comb \Selector139~0 (
	.dataa(!m_data_11),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.datae(!\active_data[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector139~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector139~0 .extended_lut = "off";
defparam \Selector139~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector139~0 .shared_arith = "off";

dffeas \active_data[12] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[12]~q ),
	.prn(vcc));
defparam \active_data[12] .is_wysiwyg = "true";
defparam \active_data[12] .power_up = "low";

cyclonev_lcell_comb \Selector138~0 (
	.dataa(!m_data_12),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.datae(!\active_data[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector138~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector138~0 .extended_lut = "off";
defparam \Selector138~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector138~0 .shared_arith = "off";

dffeas \active_data[13] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[13]~q ),
	.prn(vcc));
defparam \active_data[13] .is_wysiwyg = "true";
defparam \active_data[13] .power_up = "low";

cyclonev_lcell_comb \Selector137~0 (
	.dataa(!m_data_13),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.datae(!\active_data[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector137~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector137~0 .extended_lut = "off";
defparam \Selector137~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector137~0 .shared_arith = "off";

dffeas \active_data[14] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[14]~q ),
	.prn(vcc));
defparam \active_data[14] .is_wysiwyg = "true";
defparam \active_data[14] .power_up = "low";

cyclonev_lcell_comb \Selector136~0 (
	.dataa(!m_data_14),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.datae(!\active_data[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector136~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector136~0 .extended_lut = "off";
defparam \Selector136~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector136~0 .shared_arith = "off";

dffeas \active_data[15] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[15]~q ),
	.prn(vcc));
defparam \active_data[15] .is_wysiwyg = "true";
defparam \active_data[15] .power_up = "low";

cyclonev_lcell_comb \Selector135~0 (
	.dataa(!m_data_15),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.datae(!\active_data[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector135~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector135~0 .extended_lut = "off";
defparam \Selector135~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector135~0 .shared_arith = "off";

dffeas \active_data[16] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[16]~q ),
	.prn(vcc));
defparam \active_data[16] .is_wysiwyg = "true";
defparam \active_data[16] .power_up = "low";

cyclonev_lcell_comb \Selector134~0 (
	.dataa(!m_data_16),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.datae(!\active_data[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector134~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector134~0 .extended_lut = "off";
defparam \Selector134~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector134~0 .shared_arith = "off";

dffeas \active_data[17] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[17]~q ),
	.prn(vcc));
defparam \active_data[17] .is_wysiwyg = "true";
defparam \active_data[17] .power_up = "low";

cyclonev_lcell_comb \Selector133~0 (
	.dataa(!m_data_17),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.datae(!\active_data[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector133~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector133~0 .extended_lut = "off";
defparam \Selector133~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector133~0 .shared_arith = "off";

dffeas \active_data[18] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[18]~q ),
	.prn(vcc));
defparam \active_data[18] .is_wysiwyg = "true";
defparam \active_data[18] .power_up = "low";

cyclonev_lcell_comb \Selector132~0 (
	.dataa(!m_data_18),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.datae(!\active_data[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector132~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector132~0 .extended_lut = "off";
defparam \Selector132~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector132~0 .shared_arith = "off";

dffeas \active_data[19] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[19]~q ),
	.prn(vcc));
defparam \active_data[19] .is_wysiwyg = "true";
defparam \active_data[19] .power_up = "low";

cyclonev_lcell_comb \Selector131~0 (
	.dataa(!m_data_19),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.datae(!\active_data[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector131~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector131~0 .extended_lut = "off";
defparam \Selector131~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector131~0 .shared_arith = "off";

dffeas \active_data[20] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[20]~q ),
	.prn(vcc));
defparam \active_data[20] .is_wysiwyg = "true";
defparam \active_data[20] .power_up = "low";

cyclonev_lcell_comb \Selector130~0 (
	.dataa(!m_data_20),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.datae(!\active_data[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector130~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector130~0 .extended_lut = "off";
defparam \Selector130~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector130~0 .shared_arith = "off";

dffeas \active_data[21] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[21]~q ),
	.prn(vcc));
defparam \active_data[21] .is_wysiwyg = "true";
defparam \active_data[21] .power_up = "low";

cyclonev_lcell_comb \Selector129~0 (
	.dataa(!m_data_21),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.datae(!\active_data[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector129~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector129~0 .extended_lut = "off";
defparam \Selector129~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector129~0 .shared_arith = "off";

dffeas \active_data[22] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[22]~q ),
	.prn(vcc));
defparam \active_data[22] .is_wysiwyg = "true";
defparam \active_data[22] .power_up = "low";

cyclonev_lcell_comb \Selector128~0 (
	.dataa(!m_data_22),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.datae(!\active_data[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector128~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector128~0 .extended_lut = "off";
defparam \Selector128~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector128~0 .shared_arith = "off";

dffeas \active_data[23] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[23]~q ),
	.prn(vcc));
defparam \active_data[23] .is_wysiwyg = "true";
defparam \active_data[23] .power_up = "low";

cyclonev_lcell_comb \Selector127~0 (
	.dataa(!m_data_23),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.datae(!\active_data[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector127~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector127~0 .extended_lut = "off";
defparam \Selector127~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector127~0 .shared_arith = "off";

dffeas \active_data[24] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[24]~q ),
	.prn(vcc));
defparam \active_data[24] .is_wysiwyg = "true";
defparam \active_data[24] .power_up = "low";

cyclonev_lcell_comb \Selector126~0 (
	.dataa(!m_data_24),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.datae(!\active_data[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector126~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector126~0 .extended_lut = "off";
defparam \Selector126~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector126~0 .shared_arith = "off";

dffeas \active_data[25] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[25]~q ),
	.prn(vcc));
defparam \active_data[25] .is_wysiwyg = "true";
defparam \active_data[25] .power_up = "low";

cyclonev_lcell_comb \Selector125~0 (
	.dataa(!m_data_25),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.datae(!\active_data[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector125~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector125~0 .extended_lut = "off";
defparam \Selector125~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector125~0 .shared_arith = "off";

dffeas \active_data[26] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[26]~q ),
	.prn(vcc));
defparam \active_data[26] .is_wysiwyg = "true";
defparam \active_data[26] .power_up = "low";

cyclonev_lcell_comb \Selector124~0 (
	.dataa(!m_data_26),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.datae(!\active_data[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector124~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector124~0 .extended_lut = "off";
defparam \Selector124~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector124~0 .shared_arith = "off";

dffeas \active_data[27] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[27]~q ),
	.prn(vcc));
defparam \active_data[27] .is_wysiwyg = "true";
defparam \active_data[27] .power_up = "low";

cyclonev_lcell_comb \Selector123~0 (
	.dataa(!m_data_27),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.datae(!\active_data[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector123~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector123~0 .extended_lut = "off";
defparam \Selector123~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector123~0 .shared_arith = "off";

dffeas \active_data[28] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[28]~q ),
	.prn(vcc));
defparam \active_data[28] .is_wysiwyg = "true";
defparam \active_data[28] .power_up = "low";

cyclonev_lcell_comb \Selector122~0 (
	.dataa(!m_data_28),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.datae(!\active_data[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector122~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector122~0 .extended_lut = "off";
defparam \Selector122~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector122~0 .shared_arith = "off";

dffeas \active_data[29] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[29]~q ),
	.prn(vcc));
defparam \active_data[29] .is_wysiwyg = "true";
defparam \active_data[29] .power_up = "low";

cyclonev_lcell_comb \Selector121~0 (
	.dataa(!m_data_29),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.datae(!\active_data[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector121~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector121~0 .extended_lut = "off";
defparam \Selector121~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector121~0 .shared_arith = "off";

dffeas \active_data[30] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[30]~q ),
	.prn(vcc));
defparam \active_data[30] .is_wysiwyg = "true";
defparam \active_data[30] .power_up = "low";

cyclonev_lcell_comb \Selector120~0 (
	.dataa(!m_data_30),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.datae(!\active_data[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector120~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector120~0 .extended_lut = "off";
defparam \Selector120~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector120~0 .shared_arith = "off";

dffeas \active_data[31] (
	.clk(clk_clk),
	.d(\the_sdram_demo_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[31]~q ),
	.prn(vcc));
defparam \active_data[31] .is_wysiwyg = "true";
defparam \active_data[31] .power_up = "low";

cyclonev_lcell_comb \Selector119~0 (
	.dataa(!m_data_31),
	.datab(!\m_data[1]~0_combout ),
	.datac(!\WideOr17~0_combout ),
	.datad(!\the_sdram_demo_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.datae(!\active_data[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector119~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector119~0 .extended_lut = "off";
defparam \Selector119~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \Selector119~0 .shared_arith = "off";

endmodule

module sdram_demo_sdram_demo_sdram_input_efifo_module (
	reset_n,
	always0,
	f_pop,
	entries_1,
	entries_0,
	Equal1,
	rd_address1,
	rd_data_56,
	rd_data_57,
	entry_1_58,
	entry_0_58,
	entry_1_59,
	entry_0_59,
	entry_1_46,
	entry_0_46,
	entry_1_60,
	entry_0_60,
	entry_1_47,
	entry_0_47,
	entry_1_48,
	entry_0_48,
	entry_1_49,
	entry_0_49,
	entry_1_61,
	entry_0_61,
	entry_1_50,
	entry_0_50,
	entry_1_51,
	entry_0_51,
	entry_1_52,
	entry_0_52,
	entry_1_53,
	entry_0_53,
	entry_1_54,
	entry_0_54,
	entry_1_55,
	entry_0_55,
	Selector41,
	rd_data_36,
	rd_data_37,
	rd_data_38,
	rd_data_39,
	rd_data_40,
	rd_data_41,
	rd_data_42,
	rd_data_43,
	rd_data_44,
	rd_data_45,
	rd_data_46,
	rd_data_60,
	rd_data_32,
	rd_data_33,
	rd_data_34,
	rd_data_35,
	saved_grant_0,
	WideOr0,
	rd_data_47,
	rd_data_61,
	Equal11,
	src5_valid,
	src_valid,
	src_data_68,
	src_data_58,
	src_valid1,
	src_data_59,
	rd_data_58,
	src_data_60,
	rd_data_59,
	src_data_61,
	src_data_48,
	src_data_62,
	src_data_49,
	rd_data_48,
	src_data_50,
	rd_data_49,
	src_data_51,
	m0_write,
	rd_data_50,
	src_data_52,
	rd_data_51,
	src_data_53,
	rd_data_52,
	src_data_54,
	rd_data_53,
	src_data_55,
	rd_data_54,
	src_data_56,
	rd_data_55,
	src_data_57,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	comb,
	comb1,
	comb2,
	comb3,
	rd_data_0,
	rd_data_1,
	rd_data_2,
	rd_data_3,
	rd_data_4,
	rd_data_5,
	rd_data_6,
	rd_data_7,
	rd_data_8,
	rd_data_9,
	rd_data_10,
	rd_data_11,
	rd_data_12,
	rd_data_13,
	rd_data_14,
	rd_data_15,
	rd_data_16,
	rd_data_17,
	rd_data_18,
	rd_data_19,
	rd_data_20,
	rd_data_21,
	rd_data_22,
	rd_data_23,
	rd_data_24,
	rd_data_25,
	rd_data_26,
	rd_data_27,
	rd_data_28,
	rd_data_29,
	rd_data_30,
	rd_data_31,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	always0;
input 	f_pop;
output 	entries_1;
output 	entries_0;
output 	Equal1;
output 	rd_address1;
output 	rd_data_56;
output 	rd_data_57;
output 	entry_1_58;
output 	entry_0_58;
output 	entry_1_59;
output 	entry_0_59;
output 	entry_1_46;
output 	entry_0_46;
output 	entry_1_60;
output 	entry_0_60;
output 	entry_1_47;
output 	entry_0_47;
output 	entry_1_48;
output 	entry_0_48;
output 	entry_1_49;
output 	entry_0_49;
output 	entry_1_61;
output 	entry_0_61;
output 	entry_1_50;
output 	entry_0_50;
output 	entry_1_51;
output 	entry_0_51;
output 	entry_1_52;
output 	entry_0_52;
output 	entry_1_53;
output 	entry_0_53;
output 	entry_1_54;
output 	entry_0_54;
output 	entry_1_55;
output 	entry_0_55;
input 	Selector41;
output 	rd_data_36;
output 	rd_data_37;
output 	rd_data_38;
output 	rd_data_39;
output 	rd_data_40;
output 	rd_data_41;
output 	rd_data_42;
output 	rd_data_43;
output 	rd_data_44;
output 	rd_data_45;
output 	rd_data_46;
output 	rd_data_60;
output 	rd_data_32;
output 	rd_data_33;
output 	rd_data_34;
output 	rd_data_35;
input 	saved_grant_0;
input 	WideOr0;
output 	rd_data_47;
output 	rd_data_61;
input 	Equal11;
input 	src5_valid;
input 	src_valid;
input 	src_data_68;
input 	src_data_58;
input 	src_valid1;
input 	src_data_59;
output 	rd_data_58;
input 	src_data_60;
output 	rd_data_59;
input 	src_data_61;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
output 	rd_data_48;
input 	src_data_50;
output 	rd_data_49;
input 	src_data_51;
input 	m0_write;
output 	rd_data_50;
input 	src_data_52;
output 	rd_data_51;
input 	src_data_53;
output 	rd_data_52;
input 	src_data_54;
output 	rd_data_53;
input 	src_data_55;
output 	rd_data_54;
input 	src_data_56;
output 	rd_data_55;
input 	src_data_57;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	comb;
input 	comb1;
input 	comb2;
input 	comb3;
output 	rd_data_0;
output 	rd_data_1;
output 	rd_data_2;
output 	rd_data_3;
output 	rd_data_4;
output 	rd_data_5;
output 	rd_data_6;
output 	rd_data_7;
output 	rd_data_8;
output 	rd_data_9;
output 	rd_data_10;
output 	rd_data_11;
output 	rd_data_12;
output 	rd_data_13;
output 	rd_data_14;
output 	rd_data_15;
output 	rd_data_16;
output 	rd_data_17;
output 	rd_data_18;
output 	rd_data_19;
output 	rd_data_20;
output 	rd_data_21;
output 	rd_data_22;
output 	rd_data_23;
output 	rd_data_24;
output 	rd_data_25;
output 	rd_data_26;
output 	rd_data_27;
output 	rd_data_28;
output 	rd_data_29;
output 	rd_data_30;
output 	rd_data_31;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always2~0_combout ;
wire \always2~1_combout ;
wire \entries[1]~0_combout ;
wire \entries[0]~1_combout ;
wire \rd_address~0_combout ;
wire \wr_address~0_combout ;
wire \wr_address~q ;
wire \entry_1[61]~0_combout ;
wire \entry_1[56]~q ;
wire \entry_0[61]~0_combout ;
wire \entry_0[56]~q ;
wire \entry_1[57]~q ;
wire \entry_0[57]~q ;
wire \entry_1[36]~q ;
wire \entry_0[36]~q ;
wire \entry_1[37]~q ;
wire \entry_0[37]~q ;
wire \entry_1[38]~q ;
wire \entry_0[38]~q ;
wire \entry_1[39]~q ;
wire \entry_0[39]~q ;
wire \entry_1[40]~q ;
wire \entry_0[40]~q ;
wire \entry_1[41]~q ;
wire \entry_0[41]~q ;
wire \entry_1[42]~q ;
wire \entry_0[42]~q ;
wire \entry_1[43]~q ;
wire \entry_0[43]~q ;
wire \entry_1[44]~q ;
wire \entry_0[44]~q ;
wire \entry_1[45]~q ;
wire \entry_0[45]~q ;
wire \entry_1[32]~q ;
wire \entry_0[32]~q ;
wire \entry_1[33]~q ;
wire \entry_0[33]~q ;
wire \entry_1[34]~q ;
wire \entry_0[34]~q ;
wire \entry_1[35]~q ;
wire \entry_0[35]~q ;
wire \entry_1[0]~q ;
wire \entry_0[0]~q ;
wire \entry_1[1]~q ;
wire \entry_0[1]~q ;
wire \entry_1[2]~q ;
wire \entry_0[2]~q ;
wire \entry_1[3]~q ;
wire \entry_0[3]~q ;
wire \entry_1[4]~q ;
wire \entry_0[4]~q ;
wire \entry_1[5]~q ;
wire \entry_0[5]~q ;
wire \entry_1[6]~q ;
wire \entry_0[6]~q ;
wire \entry_1[7]~q ;
wire \entry_0[7]~q ;
wire \entry_1[8]~q ;
wire \entry_0[8]~q ;
wire \entry_1[9]~q ;
wire \entry_0[9]~q ;
wire \entry_1[10]~q ;
wire \entry_0[10]~q ;
wire \entry_1[11]~q ;
wire \entry_0[11]~q ;
wire \entry_1[12]~q ;
wire \entry_0[12]~q ;
wire \entry_1[13]~q ;
wire \entry_0[13]~q ;
wire \entry_1[14]~q ;
wire \entry_0[14]~q ;
wire \entry_1[15]~q ;
wire \entry_0[15]~q ;
wire \entry_1[16]~q ;
wire \entry_0[16]~q ;
wire \entry_1[17]~q ;
wire \entry_0[17]~q ;
wire \entry_1[18]~q ;
wire \entry_0[18]~q ;
wire \entry_1[19]~q ;
wire \entry_0[19]~q ;
wire \entry_1[20]~q ;
wire \entry_0[20]~q ;
wire \entry_1[21]~q ;
wire \entry_0[21]~q ;
wire \entry_1[22]~q ;
wire \entry_0[22]~q ;
wire \entry_1[23]~q ;
wire \entry_0[23]~q ;
wire \entry_1[24]~q ;
wire \entry_0[24]~q ;
wire \entry_1[25]~q ;
wire \entry_0[25]~q ;
wire \entry_1[26]~q ;
wire \entry_0[26]~q ;
wire \entry_1[27]~q ;
wire \entry_0[27]~q ;
wire \entry_1[28]~q ;
wire \entry_0[28]~q ;
wire \entry_1[29]~q ;
wire \entry_0[29]~q ;
wire \entry_1[30]~q ;
wire \entry_0[30]~q ;
wire \entry_1[31]~q ;
wire \entry_0[31]~q ;


dffeas \entries[1] (
	.clk(clk),
	.d(\entries[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_1),
	.prn(vcc));
defparam \entries[1] .is_wysiwyg = "true";
defparam \entries[1] .power_up = "low";

dffeas \entries[0] (
	.clk(clk),
	.d(\entries[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_0),
	.prn(vcc));
defparam \entries[0] .is_wysiwyg = "true";
defparam \entries[0] .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!entries_1),
	.datab(!entries_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal1~0 .shared_arith = "off";

dffeas rd_address(
	.clk(clk),
	.d(\rd_address~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_address1),
	.prn(vcc));
defparam rd_address.is_wysiwyg = "true";
defparam rd_address.power_up = "low";

cyclonev_lcell_comb \rd_data[56]~0 (
	.dataa(!rd_address1),
	.datab(!\entry_1[56]~q ),
	.datac(!\entry_0[56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_56),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[56]~0 .extended_lut = "off";
defparam \rd_data[56]~0 .lut_mask = 64'h2727272727272727;
defparam \rd_data[56]~0 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[57]~1 (
	.dataa(!rd_address1),
	.datab(!\entry_1[57]~q ),
	.datac(!\entry_0[57]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_57),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[57]~1 .extended_lut = "off";
defparam \rd_data[57]~1 .lut_mask = 64'h2727272727272727;
defparam \rd_data[57]~1 .shared_arith = "off";

dffeas \entry_1[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_58),
	.prn(vcc));
defparam \entry_1[58] .is_wysiwyg = "true";
defparam \entry_1[58] .power_up = "low";

dffeas \entry_0[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_58),
	.prn(vcc));
defparam \entry_0[58] .is_wysiwyg = "true";
defparam \entry_0[58] .power_up = "low";

dffeas \entry_1[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_59),
	.prn(vcc));
defparam \entry_1[59] .is_wysiwyg = "true";
defparam \entry_1[59] .power_up = "low";

dffeas \entry_0[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_59),
	.prn(vcc));
defparam \entry_0[59] .is_wysiwyg = "true";
defparam \entry_0[59] .power_up = "low";

dffeas \entry_1[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_46),
	.prn(vcc));
defparam \entry_1[46] .is_wysiwyg = "true";
defparam \entry_1[46] .power_up = "low";

dffeas \entry_0[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_46),
	.prn(vcc));
defparam \entry_0[46] .is_wysiwyg = "true";
defparam \entry_0[46] .power_up = "low";

dffeas \entry_1[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_60),
	.prn(vcc));
defparam \entry_1[60] .is_wysiwyg = "true";
defparam \entry_1[60] .power_up = "low";

dffeas \entry_0[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_60),
	.prn(vcc));
defparam \entry_0[60] .is_wysiwyg = "true";
defparam \entry_0[60] .power_up = "low";

dffeas \entry_1[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_47),
	.prn(vcc));
defparam \entry_1[47] .is_wysiwyg = "true";
defparam \entry_1[47] .power_up = "low";

dffeas \entry_0[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_47),
	.prn(vcc));
defparam \entry_0[47] .is_wysiwyg = "true";
defparam \entry_0[47] .power_up = "low";

dffeas \entry_1[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_48),
	.prn(vcc));
defparam \entry_1[48] .is_wysiwyg = "true";
defparam \entry_1[48] .power_up = "low";

dffeas \entry_0[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_48),
	.prn(vcc));
defparam \entry_0[48] .is_wysiwyg = "true";
defparam \entry_0[48] .power_up = "low";

dffeas \entry_1[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_49),
	.prn(vcc));
defparam \entry_1[49] .is_wysiwyg = "true";
defparam \entry_1[49] .power_up = "low";

dffeas \entry_0[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_49),
	.prn(vcc));
defparam \entry_0[49] .is_wysiwyg = "true";
defparam \entry_0[49] .power_up = "low";

dffeas \entry_1[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_61),
	.prn(vcc));
defparam \entry_1[61] .is_wysiwyg = "true";
defparam \entry_1[61] .power_up = "low";

dffeas \entry_0[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_61),
	.prn(vcc));
defparam \entry_0[61] .is_wysiwyg = "true";
defparam \entry_0[61] .power_up = "low";

dffeas \entry_1[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_50),
	.prn(vcc));
defparam \entry_1[50] .is_wysiwyg = "true";
defparam \entry_1[50] .power_up = "low";

dffeas \entry_0[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_50),
	.prn(vcc));
defparam \entry_0[50] .is_wysiwyg = "true";
defparam \entry_0[50] .power_up = "low";

dffeas \entry_1[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_51),
	.prn(vcc));
defparam \entry_1[51] .is_wysiwyg = "true";
defparam \entry_1[51] .power_up = "low";

dffeas \entry_0[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_51),
	.prn(vcc));
defparam \entry_0[51] .is_wysiwyg = "true";
defparam \entry_0[51] .power_up = "low";

dffeas \entry_1[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_52),
	.prn(vcc));
defparam \entry_1[52] .is_wysiwyg = "true";
defparam \entry_1[52] .power_up = "low";

dffeas \entry_0[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_52),
	.prn(vcc));
defparam \entry_0[52] .is_wysiwyg = "true";
defparam \entry_0[52] .power_up = "low";

dffeas \entry_1[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_53),
	.prn(vcc));
defparam \entry_1[53] .is_wysiwyg = "true";
defparam \entry_1[53] .power_up = "low";

dffeas \entry_0[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_53),
	.prn(vcc));
defparam \entry_0[53] .is_wysiwyg = "true";
defparam \entry_0[53] .power_up = "low";

dffeas \entry_1[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_54),
	.prn(vcc));
defparam \entry_1[54] .is_wysiwyg = "true";
defparam \entry_1[54] .power_up = "low";

dffeas \entry_0[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_54),
	.prn(vcc));
defparam \entry_0[54] .is_wysiwyg = "true";
defparam \entry_0[54] .power_up = "low";

dffeas \entry_1[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(entry_1_55),
	.prn(vcc));
defparam \entry_1[55] .is_wysiwyg = "true";
defparam \entry_1[55] .power_up = "low";

dffeas \entry_0[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(entry_0_55),
	.prn(vcc));
defparam \entry_0[55] .is_wysiwyg = "true";
defparam \entry_0[55] .power_up = "low";

cyclonev_lcell_comb \rd_data[36]~2 (
	.dataa(!rd_address1),
	.datab(!\entry_1[36]~q ),
	.datac(!\entry_0[36]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_36),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[36]~2 .extended_lut = "off";
defparam \rd_data[36]~2 .lut_mask = 64'h2727272727272727;
defparam \rd_data[36]~2 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[37]~3 (
	.dataa(!rd_address1),
	.datab(!\entry_1[37]~q ),
	.datac(!\entry_0[37]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_37),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[37]~3 .extended_lut = "off";
defparam \rd_data[37]~3 .lut_mask = 64'h2727272727272727;
defparam \rd_data[37]~3 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[38]~4 (
	.dataa(!rd_address1),
	.datab(!\entry_1[38]~q ),
	.datac(!\entry_0[38]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[38]~4 .extended_lut = "off";
defparam \rd_data[38]~4 .lut_mask = 64'h2727272727272727;
defparam \rd_data[38]~4 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[39]~5 (
	.dataa(!rd_address1),
	.datab(!\entry_1[39]~q ),
	.datac(!\entry_0[39]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[39]~5 .extended_lut = "off";
defparam \rd_data[39]~5 .lut_mask = 64'h2727272727272727;
defparam \rd_data[39]~5 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[40]~6 (
	.dataa(!rd_address1),
	.datab(!\entry_1[40]~q ),
	.datac(!\entry_0[40]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[40]~6 .extended_lut = "off";
defparam \rd_data[40]~6 .lut_mask = 64'h2727272727272727;
defparam \rd_data[40]~6 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[41]~7 (
	.dataa(!rd_address1),
	.datab(!\entry_1[41]~q ),
	.datac(!\entry_0[41]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[41]~7 .extended_lut = "off";
defparam \rd_data[41]~7 .lut_mask = 64'h2727272727272727;
defparam \rd_data[41]~7 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[42]~8 (
	.dataa(!rd_address1),
	.datab(!\entry_1[42]~q ),
	.datac(!\entry_0[42]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[42]~8 .extended_lut = "off";
defparam \rd_data[42]~8 .lut_mask = 64'h2727272727272727;
defparam \rd_data[42]~8 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[43]~9 (
	.dataa(!rd_address1),
	.datab(!\entry_1[43]~q ),
	.datac(!\entry_0[43]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[43]~9 .extended_lut = "off";
defparam \rd_data[43]~9 .lut_mask = 64'h2727272727272727;
defparam \rd_data[43]~9 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[44]~10 (
	.dataa(!rd_address1),
	.datab(!\entry_1[44]~q ),
	.datac(!\entry_0[44]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[44]~10 .extended_lut = "off";
defparam \rd_data[44]~10 .lut_mask = 64'h2727272727272727;
defparam \rd_data[44]~10 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[45]~11 (
	.dataa(!rd_address1),
	.datab(!\entry_1[45]~q ),
	.datac(!\entry_0[45]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[45]~11 .extended_lut = "off";
defparam \rd_data[45]~11 .lut_mask = 64'h2727272727272727;
defparam \rd_data[45]~11 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[46]~12 (
	.dataa(!rd_address1),
	.datab(!entry_1_46),
	.datac(!entry_0_46),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[46]~12 .extended_lut = "off";
defparam \rd_data[46]~12 .lut_mask = 64'h2727272727272727;
defparam \rd_data[46]~12 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[60]~13 (
	.dataa(!rd_address1),
	.datab(!entry_1_60),
	.datac(!entry_0_60),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_60),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[60]~13 .extended_lut = "off";
defparam \rd_data[60]~13 .lut_mask = 64'h2727272727272727;
defparam \rd_data[60]~13 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[32]~14 (
	.dataa(!rd_address1),
	.datab(!\entry_1[32]~q ),
	.datac(!\entry_0[32]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[32]~14 .extended_lut = "off";
defparam \rd_data[32]~14 .lut_mask = 64'h2727272727272727;
defparam \rd_data[32]~14 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[33]~15 (
	.dataa(!rd_address1),
	.datab(!\entry_1[33]~q ),
	.datac(!\entry_0[33]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[33]~15 .extended_lut = "off";
defparam \rd_data[33]~15 .lut_mask = 64'h2727272727272727;
defparam \rd_data[33]~15 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[34]~16 (
	.dataa(!rd_address1),
	.datab(!\entry_1[34]~q ),
	.datac(!\entry_0[34]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[34]~16 .extended_lut = "off";
defparam \rd_data[34]~16 .lut_mask = 64'h2727272727272727;
defparam \rd_data[34]~16 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[35]~17 (
	.dataa(!rd_address1),
	.datab(!\entry_1[35]~q ),
	.datac(!\entry_0[35]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[35]~17 .extended_lut = "off";
defparam \rd_data[35]~17 .lut_mask = 64'h2727272727272727;
defparam \rd_data[35]~17 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[47]~18 (
	.dataa(!rd_address1),
	.datab(!entry_1_47),
	.datac(!entry_0_47),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[47]~18 .extended_lut = "off";
defparam \rd_data[47]~18 .lut_mask = 64'h2727272727272727;
defparam \rd_data[47]~18 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[61]~19 (
	.dataa(!rd_address1),
	.datab(!entry_1_61),
	.datac(!entry_0_61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_61),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[61]~19 .extended_lut = "off";
defparam \rd_data[61]~19 .lut_mask = 64'h2727272727272727;
defparam \rd_data[61]~19 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[58]~20 (
	.dataa(!rd_address1),
	.datab(!entry_1_58),
	.datac(!entry_0_58),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_58),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[58]~20 .extended_lut = "off";
defparam \rd_data[58]~20 .lut_mask = 64'h2727272727272727;
defparam \rd_data[58]~20 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[59]~21 (
	.dataa(!rd_address1),
	.datab(!entry_1_59),
	.datac(!entry_0_59),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_59),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[59]~21 .extended_lut = "off";
defparam \rd_data[59]~21 .lut_mask = 64'h2727272727272727;
defparam \rd_data[59]~21 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[48]~22 (
	.dataa(!rd_address1),
	.datab(!entry_1_48),
	.datac(!entry_0_48),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[48]~22 .extended_lut = "off";
defparam \rd_data[48]~22 .lut_mask = 64'h2727272727272727;
defparam \rd_data[48]~22 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[49]~23 (
	.dataa(!rd_address1),
	.datab(!entry_1_49),
	.datac(!entry_0_49),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[49]~23 .extended_lut = "off";
defparam \rd_data[49]~23 .lut_mask = 64'h2727272727272727;
defparam \rd_data[49]~23 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[50]~24 (
	.dataa(!rd_address1),
	.datab(!entry_1_50),
	.datac(!entry_0_50),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[50]~24 .extended_lut = "off";
defparam \rd_data[50]~24 .lut_mask = 64'h2727272727272727;
defparam \rd_data[50]~24 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[51]~25 (
	.dataa(!rd_address1),
	.datab(!entry_1_51),
	.datac(!entry_0_51),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[51]~25 .extended_lut = "off";
defparam \rd_data[51]~25 .lut_mask = 64'h2727272727272727;
defparam \rd_data[51]~25 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[52]~26 (
	.dataa(!rd_address1),
	.datab(!entry_1_52),
	.datac(!entry_0_52),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_52),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[52]~26 .extended_lut = "off";
defparam \rd_data[52]~26 .lut_mask = 64'h2727272727272727;
defparam \rd_data[52]~26 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[53]~27 (
	.dataa(!rd_address1),
	.datab(!entry_1_53),
	.datac(!entry_0_53),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_53),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[53]~27 .extended_lut = "off";
defparam \rd_data[53]~27 .lut_mask = 64'h2727272727272727;
defparam \rd_data[53]~27 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[54]~28 (
	.dataa(!rd_address1),
	.datab(!entry_1_54),
	.datac(!entry_0_54),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_54),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[54]~28 .extended_lut = "off";
defparam \rd_data[54]~28 .lut_mask = 64'h2727272727272727;
defparam \rd_data[54]~28 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[55]~29 (
	.dataa(!rd_address1),
	.datab(!entry_1_55),
	.datac(!entry_0_55),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_55),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[55]~29 .extended_lut = "off";
defparam \rd_data[55]~29 .lut_mask = 64'h2727272727272727;
defparam \rd_data[55]~29 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[0]~30 (
	.dataa(!rd_address1),
	.datab(!\entry_1[0]~q ),
	.datac(!\entry_0[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[0]~30 .extended_lut = "off";
defparam \rd_data[0]~30 .lut_mask = 64'h2727272727272727;
defparam \rd_data[0]~30 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[1]~31 (
	.dataa(!rd_address1),
	.datab(!\entry_1[1]~q ),
	.datac(!\entry_0[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[1]~31 .extended_lut = "off";
defparam \rd_data[1]~31 .lut_mask = 64'h2727272727272727;
defparam \rd_data[1]~31 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[2]~32 (
	.dataa(!rd_address1),
	.datab(!\entry_1[2]~q ),
	.datac(!\entry_0[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[2]~32 .extended_lut = "off";
defparam \rd_data[2]~32 .lut_mask = 64'h2727272727272727;
defparam \rd_data[2]~32 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[3]~33 (
	.dataa(!rd_address1),
	.datab(!\entry_1[3]~q ),
	.datac(!\entry_0[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[3]~33 .extended_lut = "off";
defparam \rd_data[3]~33 .lut_mask = 64'h2727272727272727;
defparam \rd_data[3]~33 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[4]~34 (
	.dataa(!rd_address1),
	.datab(!\entry_1[4]~q ),
	.datac(!\entry_0[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[4]~34 .extended_lut = "off";
defparam \rd_data[4]~34 .lut_mask = 64'h2727272727272727;
defparam \rd_data[4]~34 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[5]~35 (
	.dataa(!rd_address1),
	.datab(!\entry_1[5]~q ),
	.datac(!\entry_0[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[5]~35 .extended_lut = "off";
defparam \rd_data[5]~35 .lut_mask = 64'h2727272727272727;
defparam \rd_data[5]~35 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[6]~36 (
	.dataa(!rd_address1),
	.datab(!\entry_1[6]~q ),
	.datac(!\entry_0[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[6]~36 .extended_lut = "off";
defparam \rd_data[6]~36 .lut_mask = 64'h2727272727272727;
defparam \rd_data[6]~36 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[7]~37 (
	.dataa(!rd_address1),
	.datab(!\entry_1[7]~q ),
	.datac(!\entry_0[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[7]~37 .extended_lut = "off";
defparam \rd_data[7]~37 .lut_mask = 64'h2727272727272727;
defparam \rd_data[7]~37 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[8]~38 (
	.dataa(!rd_address1),
	.datab(!\entry_1[8]~q ),
	.datac(!\entry_0[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[8]~38 .extended_lut = "off";
defparam \rd_data[8]~38 .lut_mask = 64'h2727272727272727;
defparam \rd_data[8]~38 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[9]~39 (
	.dataa(!rd_address1),
	.datab(!\entry_1[9]~q ),
	.datac(!\entry_0[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[9]~39 .extended_lut = "off";
defparam \rd_data[9]~39 .lut_mask = 64'h2727272727272727;
defparam \rd_data[9]~39 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[10]~40 (
	.dataa(!rd_address1),
	.datab(!\entry_1[10]~q ),
	.datac(!\entry_0[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[10]~40 .extended_lut = "off";
defparam \rd_data[10]~40 .lut_mask = 64'h2727272727272727;
defparam \rd_data[10]~40 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[11]~41 (
	.dataa(!rd_address1),
	.datab(!\entry_1[11]~q ),
	.datac(!\entry_0[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[11]~41 .extended_lut = "off";
defparam \rd_data[11]~41 .lut_mask = 64'h2727272727272727;
defparam \rd_data[11]~41 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[12]~42 (
	.dataa(!rd_address1),
	.datab(!\entry_1[12]~q ),
	.datac(!\entry_0[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[12]~42 .extended_lut = "off";
defparam \rd_data[12]~42 .lut_mask = 64'h2727272727272727;
defparam \rd_data[12]~42 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[13]~43 (
	.dataa(!rd_address1),
	.datab(!\entry_1[13]~q ),
	.datac(!\entry_0[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[13]~43 .extended_lut = "off";
defparam \rd_data[13]~43 .lut_mask = 64'h2727272727272727;
defparam \rd_data[13]~43 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[14]~44 (
	.dataa(!rd_address1),
	.datab(!\entry_1[14]~q ),
	.datac(!\entry_0[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[14]~44 .extended_lut = "off";
defparam \rd_data[14]~44 .lut_mask = 64'h2727272727272727;
defparam \rd_data[14]~44 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[15]~45 (
	.dataa(!rd_address1),
	.datab(!\entry_1[15]~q ),
	.datac(!\entry_0[15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[15]~45 .extended_lut = "off";
defparam \rd_data[15]~45 .lut_mask = 64'h2727272727272727;
defparam \rd_data[15]~45 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[16]~46 (
	.dataa(!rd_address1),
	.datab(!\entry_1[16]~q ),
	.datac(!\entry_0[16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[16]~46 .extended_lut = "off";
defparam \rd_data[16]~46 .lut_mask = 64'h2727272727272727;
defparam \rd_data[16]~46 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[17]~47 (
	.dataa(!rd_address1),
	.datab(!\entry_1[17]~q ),
	.datac(!\entry_0[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[17]~47 .extended_lut = "off";
defparam \rd_data[17]~47 .lut_mask = 64'h2727272727272727;
defparam \rd_data[17]~47 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[18]~48 (
	.dataa(!rd_address1),
	.datab(!\entry_1[18]~q ),
	.datac(!\entry_0[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[18]~48 .extended_lut = "off";
defparam \rd_data[18]~48 .lut_mask = 64'h2727272727272727;
defparam \rd_data[18]~48 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[19]~49 (
	.dataa(!rd_address1),
	.datab(!\entry_1[19]~q ),
	.datac(!\entry_0[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[19]~49 .extended_lut = "off";
defparam \rd_data[19]~49 .lut_mask = 64'h2727272727272727;
defparam \rd_data[19]~49 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[20]~50 (
	.dataa(!rd_address1),
	.datab(!\entry_1[20]~q ),
	.datac(!\entry_0[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[20]~50 .extended_lut = "off";
defparam \rd_data[20]~50 .lut_mask = 64'h2727272727272727;
defparam \rd_data[20]~50 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[21]~51 (
	.dataa(!rd_address1),
	.datab(!\entry_1[21]~q ),
	.datac(!\entry_0[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[21]~51 .extended_lut = "off";
defparam \rd_data[21]~51 .lut_mask = 64'h2727272727272727;
defparam \rd_data[21]~51 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[22]~52 (
	.dataa(!rd_address1),
	.datab(!\entry_1[22]~q ),
	.datac(!\entry_0[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[22]~52 .extended_lut = "off";
defparam \rd_data[22]~52 .lut_mask = 64'h2727272727272727;
defparam \rd_data[22]~52 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[23]~53 (
	.dataa(!rd_address1),
	.datab(!\entry_1[23]~q ),
	.datac(!\entry_0[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[23]~53 .extended_lut = "off";
defparam \rd_data[23]~53 .lut_mask = 64'h2727272727272727;
defparam \rd_data[23]~53 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[24]~54 (
	.dataa(!rd_address1),
	.datab(!\entry_1[24]~q ),
	.datac(!\entry_0[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[24]~54 .extended_lut = "off";
defparam \rd_data[24]~54 .lut_mask = 64'h2727272727272727;
defparam \rd_data[24]~54 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[25]~55 (
	.dataa(!rd_address1),
	.datab(!\entry_1[25]~q ),
	.datac(!\entry_0[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[25]~55 .extended_lut = "off";
defparam \rd_data[25]~55 .lut_mask = 64'h2727272727272727;
defparam \rd_data[25]~55 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[26]~56 (
	.dataa(!rd_address1),
	.datab(!\entry_1[26]~q ),
	.datac(!\entry_0[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[26]~56 .extended_lut = "off";
defparam \rd_data[26]~56 .lut_mask = 64'h2727272727272727;
defparam \rd_data[26]~56 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[27]~57 (
	.dataa(!rd_address1),
	.datab(!\entry_1[27]~q ),
	.datac(!\entry_0[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[27]~57 .extended_lut = "off";
defparam \rd_data[27]~57 .lut_mask = 64'h2727272727272727;
defparam \rd_data[27]~57 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[28]~58 (
	.dataa(!rd_address1),
	.datab(!\entry_1[28]~q ),
	.datac(!\entry_0[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[28]~58 .extended_lut = "off";
defparam \rd_data[28]~58 .lut_mask = 64'h2727272727272727;
defparam \rd_data[28]~58 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[29]~59 (
	.dataa(!rd_address1),
	.datab(!\entry_1[29]~q ),
	.datac(!\entry_0[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[29]~59 .extended_lut = "off";
defparam \rd_data[29]~59 .lut_mask = 64'h2727272727272727;
defparam \rd_data[29]~59 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[30]~60 (
	.dataa(!rd_address1),
	.datab(!\entry_1[30]~q ),
	.datac(!\entry_0[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[30]~60 .extended_lut = "off";
defparam \rd_data[30]~60 .lut_mask = 64'h2727272727272727;
defparam \rd_data[30]~60 .shared_arith = "off";

cyclonev_lcell_comb \rd_data[31]~61 (
	.dataa(!rd_address1),
	.datab(!\entry_1[31]~q ),
	.datac(!\entry_0[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rd_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_data[31]~61 .extended_lut = "off";
defparam \rd_data[31]~61 .lut_mask = 64'h2727272727272727;
defparam \rd_data[31]~61 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!always0),
	.datab(!saved_grant_0),
	.datac(!src_data_68),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~1 (
	.dataa(!saved_grant_0),
	.datab(!WideOr0),
	.datac(!Equal11),
	.datad(!src5_valid),
	.datae(!src_valid),
	.dataf(!\always2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'hFFFFFFFFF7FFFFFF;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \entries[1]~0 (
	.dataa(!f_pop),
	.datab(!entries_1),
	.datac(!entries_0),
	.datad(!Selector41),
	.datae(!\always2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\entries[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \entries[1]~0 .extended_lut = "off";
defparam \entries[1]~0 .lut_mask = 64'h9669699696696996;
defparam \entries[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \entries[0]~1 (
	.dataa(!f_pop),
	.datab(!entries_0),
	.datac(!Selector41),
	.datad(!\always2~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\entries[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \entries[0]~1 .extended_lut = "off";
defparam \entries[0]~1 .lut_mask = 64'h6996699669966996;
defparam \entries[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \rd_address~0 (
	.dataa(!f_pop),
	.datab(!rd_address1),
	.datac(!Selector41),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_address~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_address~0 .extended_lut = "off";
defparam \rd_address~0 .lut_mask = 64'h9696969696969696;
defparam \rd_address~0 .shared_arith = "off";

cyclonev_lcell_comb \wr_address~0 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!\wr_address~q ),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_address~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_address~0 .extended_lut = "off";
defparam \wr_address~0 .lut_mask = 64'h9669699696696996;
defparam \wr_address~0 .shared_arith = "off";

dffeas wr_address(
	.clk(clk),
	.d(\wr_address~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_address~q ),
	.prn(vcc));
defparam wr_address.is_wysiwyg = "true";
defparam wr_address.power_up = "low";

cyclonev_lcell_comb \entry_1[61]~0 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!\wr_address~q ),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\entry_1[61]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \entry_1[61]~0 .extended_lut = "off";
defparam \entry_1[61]~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \entry_1[61]~0 .shared_arith = "off";

dffeas \entry_1[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[56]~q ),
	.prn(vcc));
defparam \entry_1[56] .is_wysiwyg = "true";
defparam \entry_1[56] .power_up = "low";

cyclonev_lcell_comb \entry_0[61]~0 (
	.dataa(!WideOr0),
	.datab(!src_valid1),
	.datac(!src_valid),
	.datad(!\wr_address~q ),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\entry_0[61]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \entry_0[61]~0 .extended_lut = "off";
defparam \entry_0[61]~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \entry_0[61]~0 .shared_arith = "off";

dffeas \entry_0[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[56]~q ),
	.prn(vcc));
defparam \entry_0[56] .is_wysiwyg = "true";
defparam \entry_0[56] .power_up = "low";

dffeas \entry_1[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[57]~q ),
	.prn(vcc));
defparam \entry_1[57] .is_wysiwyg = "true";
defparam \entry_1[57] .power_up = "low";

dffeas \entry_0[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[57]~q ),
	.prn(vcc));
defparam \entry_0[57] .is_wysiwyg = "true";
defparam \entry_0[57] .power_up = "low";

dffeas \entry_1[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[36]~q ),
	.prn(vcc));
defparam \entry_1[36] .is_wysiwyg = "true";
defparam \entry_1[36] .power_up = "low";

dffeas \entry_0[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[36]~q ),
	.prn(vcc));
defparam \entry_0[36] .is_wysiwyg = "true";
defparam \entry_0[36] .power_up = "low";

dffeas \entry_1[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[37]~q ),
	.prn(vcc));
defparam \entry_1[37] .is_wysiwyg = "true";
defparam \entry_1[37] .power_up = "low";

dffeas \entry_0[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[37]~q ),
	.prn(vcc));
defparam \entry_0[37] .is_wysiwyg = "true";
defparam \entry_0[37] .power_up = "low";

dffeas \entry_1[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[38]~q ),
	.prn(vcc));
defparam \entry_1[38] .is_wysiwyg = "true";
defparam \entry_1[38] .power_up = "low";

dffeas \entry_0[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[38]~q ),
	.prn(vcc));
defparam \entry_0[38] .is_wysiwyg = "true";
defparam \entry_0[38] .power_up = "low";

dffeas \entry_1[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[39]~q ),
	.prn(vcc));
defparam \entry_1[39] .is_wysiwyg = "true";
defparam \entry_1[39] .power_up = "low";

dffeas \entry_0[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[39]~q ),
	.prn(vcc));
defparam \entry_0[39] .is_wysiwyg = "true";
defparam \entry_0[39] .power_up = "low";

dffeas \entry_1[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[40]~q ),
	.prn(vcc));
defparam \entry_1[40] .is_wysiwyg = "true";
defparam \entry_1[40] .power_up = "low";

dffeas \entry_0[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[40]~q ),
	.prn(vcc));
defparam \entry_0[40] .is_wysiwyg = "true";
defparam \entry_0[40] .power_up = "low";

dffeas \entry_1[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[41]~q ),
	.prn(vcc));
defparam \entry_1[41] .is_wysiwyg = "true";
defparam \entry_1[41] .power_up = "low";

dffeas \entry_0[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[41]~q ),
	.prn(vcc));
defparam \entry_0[41] .is_wysiwyg = "true";
defparam \entry_0[41] .power_up = "low";

dffeas \entry_1[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[42]~q ),
	.prn(vcc));
defparam \entry_1[42] .is_wysiwyg = "true";
defparam \entry_1[42] .power_up = "low";

dffeas \entry_0[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[42]~q ),
	.prn(vcc));
defparam \entry_0[42] .is_wysiwyg = "true";
defparam \entry_0[42] .power_up = "low";

dffeas \entry_1[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[43]~q ),
	.prn(vcc));
defparam \entry_1[43] .is_wysiwyg = "true";
defparam \entry_1[43] .power_up = "low";

dffeas \entry_0[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[43]~q ),
	.prn(vcc));
defparam \entry_0[43] .is_wysiwyg = "true";
defparam \entry_0[43] .power_up = "low";

dffeas \entry_1[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[44]~q ),
	.prn(vcc));
defparam \entry_1[44] .is_wysiwyg = "true";
defparam \entry_1[44] .power_up = "low";

dffeas \entry_0[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[44]~q ),
	.prn(vcc));
defparam \entry_0[44] .is_wysiwyg = "true";
defparam \entry_0[44] .power_up = "low";

dffeas \entry_1[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[45]~q ),
	.prn(vcc));
defparam \entry_1[45] .is_wysiwyg = "true";
defparam \entry_1[45] .power_up = "low";

dffeas \entry_0[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[45]~q ),
	.prn(vcc));
defparam \entry_0[45] .is_wysiwyg = "true";
defparam \entry_0[45] .power_up = "low";

dffeas \entry_1[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[32]~q ),
	.prn(vcc));
defparam \entry_1[32] .is_wysiwyg = "true";
defparam \entry_1[32] .power_up = "low";

dffeas \entry_0[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[32]~q ),
	.prn(vcc));
defparam \entry_0[32] .is_wysiwyg = "true";
defparam \entry_0[32] .power_up = "low";

dffeas \entry_1[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[33]~q ),
	.prn(vcc));
defparam \entry_1[33] .is_wysiwyg = "true";
defparam \entry_1[33] .power_up = "low";

dffeas \entry_0[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[33]~q ),
	.prn(vcc));
defparam \entry_0[33] .is_wysiwyg = "true";
defparam \entry_0[33] .power_up = "low";

dffeas \entry_1[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[34]~q ),
	.prn(vcc));
defparam \entry_1[34] .is_wysiwyg = "true";
defparam \entry_1[34] .power_up = "low";

dffeas \entry_0[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[34]~q ),
	.prn(vcc));
defparam \entry_0[34] .is_wysiwyg = "true";
defparam \entry_0[34] .power_up = "low";

dffeas \entry_1[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[35]~q ),
	.prn(vcc));
defparam \entry_1[35] .is_wysiwyg = "true";
defparam \entry_1[35] .power_up = "low";

dffeas \entry_0[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[35]~q ),
	.prn(vcc));
defparam \entry_0[35] .is_wysiwyg = "true";
defparam \entry_0[35] .power_up = "low";

dffeas \entry_1[0] (
	.clk(clk),
	.d(src_payload),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[0]~q ),
	.prn(vcc));
defparam \entry_1[0] .is_wysiwyg = "true";
defparam \entry_1[0] .power_up = "low";

dffeas \entry_0[0] (
	.clk(clk),
	.d(src_payload),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[0]~q ),
	.prn(vcc));
defparam \entry_0[0] .is_wysiwyg = "true";
defparam \entry_0[0] .power_up = "low";

dffeas \entry_1[1] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[1]~q ),
	.prn(vcc));
defparam \entry_1[1] .is_wysiwyg = "true";
defparam \entry_1[1] .power_up = "low";

dffeas \entry_0[1] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[1]~q ),
	.prn(vcc));
defparam \entry_0[1] .is_wysiwyg = "true";
defparam \entry_0[1] .power_up = "low";

dffeas \entry_1[2] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[2]~q ),
	.prn(vcc));
defparam \entry_1[2] .is_wysiwyg = "true";
defparam \entry_1[2] .power_up = "low";

dffeas \entry_0[2] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[2]~q ),
	.prn(vcc));
defparam \entry_0[2] .is_wysiwyg = "true";
defparam \entry_0[2] .power_up = "low";

dffeas \entry_1[3] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[3]~q ),
	.prn(vcc));
defparam \entry_1[3] .is_wysiwyg = "true";
defparam \entry_1[3] .power_up = "low";

dffeas \entry_0[3] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[3]~q ),
	.prn(vcc));
defparam \entry_0[3] .is_wysiwyg = "true";
defparam \entry_0[3] .power_up = "low";

dffeas \entry_1[4] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[4]~q ),
	.prn(vcc));
defparam \entry_1[4] .is_wysiwyg = "true";
defparam \entry_1[4] .power_up = "low";

dffeas \entry_0[4] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[4]~q ),
	.prn(vcc));
defparam \entry_0[4] .is_wysiwyg = "true";
defparam \entry_0[4] .power_up = "low";

dffeas \entry_1[5] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[5]~q ),
	.prn(vcc));
defparam \entry_1[5] .is_wysiwyg = "true";
defparam \entry_1[5] .power_up = "low";

dffeas \entry_0[5] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[5]~q ),
	.prn(vcc));
defparam \entry_0[5] .is_wysiwyg = "true";
defparam \entry_0[5] .power_up = "low";

dffeas \entry_1[6] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[6]~q ),
	.prn(vcc));
defparam \entry_1[6] .is_wysiwyg = "true";
defparam \entry_1[6] .power_up = "low";

dffeas \entry_0[6] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[6]~q ),
	.prn(vcc));
defparam \entry_0[6] .is_wysiwyg = "true";
defparam \entry_0[6] .power_up = "low";

dffeas \entry_1[7] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[7]~q ),
	.prn(vcc));
defparam \entry_1[7] .is_wysiwyg = "true";
defparam \entry_1[7] .power_up = "low";

dffeas \entry_0[7] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[7]~q ),
	.prn(vcc));
defparam \entry_0[7] .is_wysiwyg = "true";
defparam \entry_0[7] .power_up = "low";

dffeas \entry_1[8] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[8]~q ),
	.prn(vcc));
defparam \entry_1[8] .is_wysiwyg = "true";
defparam \entry_1[8] .power_up = "low";

dffeas \entry_0[8] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[8]~q ),
	.prn(vcc));
defparam \entry_0[8] .is_wysiwyg = "true";
defparam \entry_0[8] .power_up = "low";

dffeas \entry_1[9] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[9]~q ),
	.prn(vcc));
defparam \entry_1[9] .is_wysiwyg = "true";
defparam \entry_1[9] .power_up = "low";

dffeas \entry_0[9] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[9]~q ),
	.prn(vcc));
defparam \entry_0[9] .is_wysiwyg = "true";
defparam \entry_0[9] .power_up = "low";

dffeas \entry_1[10] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[10]~q ),
	.prn(vcc));
defparam \entry_1[10] .is_wysiwyg = "true";
defparam \entry_1[10] .power_up = "low";

dffeas \entry_0[10] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[10]~q ),
	.prn(vcc));
defparam \entry_0[10] .is_wysiwyg = "true";
defparam \entry_0[10] .power_up = "low";

dffeas \entry_1[11] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[11]~q ),
	.prn(vcc));
defparam \entry_1[11] .is_wysiwyg = "true";
defparam \entry_1[11] .power_up = "low";

dffeas \entry_0[11] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[11]~q ),
	.prn(vcc));
defparam \entry_0[11] .is_wysiwyg = "true";
defparam \entry_0[11] .power_up = "low";

dffeas \entry_1[12] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[12]~q ),
	.prn(vcc));
defparam \entry_1[12] .is_wysiwyg = "true";
defparam \entry_1[12] .power_up = "low";

dffeas \entry_0[12] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[12]~q ),
	.prn(vcc));
defparam \entry_0[12] .is_wysiwyg = "true";
defparam \entry_0[12] .power_up = "low";

dffeas \entry_1[13] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[13]~q ),
	.prn(vcc));
defparam \entry_1[13] .is_wysiwyg = "true";
defparam \entry_1[13] .power_up = "low";

dffeas \entry_0[13] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[13]~q ),
	.prn(vcc));
defparam \entry_0[13] .is_wysiwyg = "true";
defparam \entry_0[13] .power_up = "low";

dffeas \entry_1[14] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[14]~q ),
	.prn(vcc));
defparam \entry_1[14] .is_wysiwyg = "true";
defparam \entry_1[14] .power_up = "low";

dffeas \entry_0[14] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[14]~q ),
	.prn(vcc));
defparam \entry_0[14] .is_wysiwyg = "true";
defparam \entry_0[14] .power_up = "low";

dffeas \entry_1[15] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[15]~q ),
	.prn(vcc));
defparam \entry_1[15] .is_wysiwyg = "true";
defparam \entry_1[15] .power_up = "low";

dffeas \entry_0[15] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[15]~q ),
	.prn(vcc));
defparam \entry_0[15] .is_wysiwyg = "true";
defparam \entry_0[15] .power_up = "low";

dffeas \entry_1[16] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[16]~q ),
	.prn(vcc));
defparam \entry_1[16] .is_wysiwyg = "true";
defparam \entry_1[16] .power_up = "low";

dffeas \entry_0[16] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[16]~q ),
	.prn(vcc));
defparam \entry_0[16] .is_wysiwyg = "true";
defparam \entry_0[16] .power_up = "low";

dffeas \entry_1[17] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[17]~q ),
	.prn(vcc));
defparam \entry_1[17] .is_wysiwyg = "true";
defparam \entry_1[17] .power_up = "low";

dffeas \entry_0[17] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[17]~q ),
	.prn(vcc));
defparam \entry_0[17] .is_wysiwyg = "true";
defparam \entry_0[17] .power_up = "low";

dffeas \entry_1[18] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[18]~q ),
	.prn(vcc));
defparam \entry_1[18] .is_wysiwyg = "true";
defparam \entry_1[18] .power_up = "low";

dffeas \entry_0[18] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[18]~q ),
	.prn(vcc));
defparam \entry_0[18] .is_wysiwyg = "true";
defparam \entry_0[18] .power_up = "low";

dffeas \entry_1[19] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[19]~q ),
	.prn(vcc));
defparam \entry_1[19] .is_wysiwyg = "true";
defparam \entry_1[19] .power_up = "low";

dffeas \entry_0[19] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[19]~q ),
	.prn(vcc));
defparam \entry_0[19] .is_wysiwyg = "true";
defparam \entry_0[19] .power_up = "low";

dffeas \entry_1[20] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[20]~q ),
	.prn(vcc));
defparam \entry_1[20] .is_wysiwyg = "true";
defparam \entry_1[20] .power_up = "low";

dffeas \entry_0[20] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[20]~q ),
	.prn(vcc));
defparam \entry_0[20] .is_wysiwyg = "true";
defparam \entry_0[20] .power_up = "low";

dffeas \entry_1[21] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[21]~q ),
	.prn(vcc));
defparam \entry_1[21] .is_wysiwyg = "true";
defparam \entry_1[21] .power_up = "low";

dffeas \entry_0[21] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[21]~q ),
	.prn(vcc));
defparam \entry_0[21] .is_wysiwyg = "true";
defparam \entry_0[21] .power_up = "low";

dffeas \entry_1[22] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[22]~q ),
	.prn(vcc));
defparam \entry_1[22] .is_wysiwyg = "true";
defparam \entry_1[22] .power_up = "low";

dffeas \entry_0[22] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[22]~q ),
	.prn(vcc));
defparam \entry_0[22] .is_wysiwyg = "true";
defparam \entry_0[22] .power_up = "low";

dffeas \entry_1[23] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[23]~q ),
	.prn(vcc));
defparam \entry_1[23] .is_wysiwyg = "true";
defparam \entry_1[23] .power_up = "low";

dffeas \entry_0[23] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[23]~q ),
	.prn(vcc));
defparam \entry_0[23] .is_wysiwyg = "true";
defparam \entry_0[23] .power_up = "low";

dffeas \entry_1[24] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[24]~q ),
	.prn(vcc));
defparam \entry_1[24] .is_wysiwyg = "true";
defparam \entry_1[24] .power_up = "low";

dffeas \entry_0[24] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[24]~q ),
	.prn(vcc));
defparam \entry_0[24] .is_wysiwyg = "true";
defparam \entry_0[24] .power_up = "low";

dffeas \entry_1[25] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[25]~q ),
	.prn(vcc));
defparam \entry_1[25] .is_wysiwyg = "true";
defparam \entry_1[25] .power_up = "low";

dffeas \entry_0[25] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[25]~q ),
	.prn(vcc));
defparam \entry_0[25] .is_wysiwyg = "true";
defparam \entry_0[25] .power_up = "low";

dffeas \entry_1[26] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[26]~q ),
	.prn(vcc));
defparam \entry_1[26] .is_wysiwyg = "true";
defparam \entry_1[26] .power_up = "low";

dffeas \entry_0[26] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[26]~q ),
	.prn(vcc));
defparam \entry_0[26] .is_wysiwyg = "true";
defparam \entry_0[26] .power_up = "low";

dffeas \entry_1[27] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[27]~q ),
	.prn(vcc));
defparam \entry_1[27] .is_wysiwyg = "true";
defparam \entry_1[27] .power_up = "low";

dffeas \entry_0[27] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[27]~q ),
	.prn(vcc));
defparam \entry_0[27] .is_wysiwyg = "true";
defparam \entry_0[27] .power_up = "low";

dffeas \entry_1[28] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[28]~q ),
	.prn(vcc));
defparam \entry_1[28] .is_wysiwyg = "true";
defparam \entry_1[28] .power_up = "low";

dffeas \entry_0[28] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[28]~q ),
	.prn(vcc));
defparam \entry_0[28] .is_wysiwyg = "true";
defparam \entry_0[28] .power_up = "low";

dffeas \entry_1[29] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[29]~q ),
	.prn(vcc));
defparam \entry_1[29] .is_wysiwyg = "true";
defparam \entry_1[29] .power_up = "low";

dffeas \entry_0[29] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[29]~q ),
	.prn(vcc));
defparam \entry_0[29] .is_wysiwyg = "true";
defparam \entry_0[29] .power_up = "low";

dffeas \entry_1[30] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[30]~q ),
	.prn(vcc));
defparam \entry_1[30] .is_wysiwyg = "true";
defparam \entry_1[30] .power_up = "low";

dffeas \entry_0[30] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[30]~q ),
	.prn(vcc));
defparam \entry_0[30] .is_wysiwyg = "true";
defparam \entry_0[30] .power_up = "low";

dffeas \entry_1[31] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[31]~q ),
	.prn(vcc));
defparam \entry_1[31] .is_wysiwyg = "true";
defparam \entry_1[31] .power_up = "low";

dffeas \entry_0[31] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[31]~q ),
	.prn(vcc));
defparam \entry_0[31] .is_wysiwyg = "true";
defparam \entry_0[31] .power_up = "low";

endmodule

module sdram_demo_sdram_demo_sw (
	W_alu_result_2,
	W_alu_result_3,
	r_sync_rst,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk_clk,
	sw_export_0,
	sw_export_1,
	sw_export_2,
	sw_export_3,
	sw_export_4,
	sw_export_5,
	sw_export_6,
	sw_export_7)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	r_sync_rst;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk_clk;
input 	sw_export_0;
input 	sw_export_1;
input 	sw_export_2;
input 	sw_export_3;
input 	sw_export_4;
input 	sw_export_5;
input 	sw_export_6;
input 	sw_export_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!W_alu_result_2),
	.datab(!W_alu_result_3),
	.datac(!sw_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[7] .shared_arith = "off";

endmodule
