-- tb: glitch01
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_GLITCHY IS
END TB_GLITCHY;

ARCHITECTURE TB OF TB_GLITCHY IS
    SIGNAL IN0 : STD_LOGIC := '0';
    SIGNAL IN1 : STD_LOGIC := '0';
    SIGNAL SEL : STD_LOGIC := '0';
    SIGNAL Z : STD_LOGIC := '0';
    SIGNAL Z_EXPECT : STD_LOGIC := '0';

    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    GLITCHY_UNIT : ENTITY WORK.GLITCHY
        PORT MAP (IN0 => IN0, IN1 => IN1, SEL => SEL, Z => Z);

    PROCESS
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE GOOD_NUM : BOOLEAN;
        VARIABLE SEPARATOR : CHARACTER;

        VARIABLE INPUT_IN0 : STD_LOGIC;
        VARIABLE INPUT_IN1 : STD_LOGIC;
        VARIABLE INPUT_SEL : STD_LOGIC;
        VARIABLE INPUT_Z : STD_LOGIC;
    BEGIN
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("SEL,IN0,IN1,Z,Z_EXPECT"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_SEL, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; -- header

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_IN0, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT("FAILED! invalid assignment for IN1");

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_IN1);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_Z);

            SEL <= INPUT_SEL;
            IN0 <= INPUT_IN0;
            IN1 <= INPUT_IN1;
            Z_EXPECT <= INPUT_Z;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, SEL);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, IN0);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, IN1);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, Z);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, Z_EXPECT);
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);
        END LOOP;
        FILE_CLOSE(OUTPUT_BUF);
        FILE_CLOSE(INPUT_BUF);
        WAIT;
    END PROCESS;
END TB;
