-- hw adaptation for DE1SoC board (cycloneV)
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DE1SOC_SHIFTER IS
PORT( SW_D : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
    ; KEY_C : IN STD_LOGIC
    ; LED_S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END DE1SOC_SHIFTER;

ARCHITECTURE DE1SOC OF DE1SOC_SHIFTER IS
    SIGNAL D : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL C : STD_LOGIC;
    SIGNAL S : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

    SHIFTER_UNIT : ENTITY WORK.SHIFTER
        PORT MAP (D => D, C => C, S => S);

    -- IN
    D <= SW_D;
    C <= NOT KEY_C;

    -- OUT
    LED_S <= S;
END DE1SOC;
