// ported from a DE2-115 demo
//
// Implements the augmented Nios II system for the DE2-115 board.
// Inputs:SW7−0 are parallel port inputs to the Nios II system.
//        CLOCK_50 is the system clock.
//        KEY0 is the active-low system reset.
// Outputs:   LEDG7−0 are parallel port outputs from the Nios II system.
//        SDRAM ports correspond to the signals in Figure 2; their names are those
//        used in the DE2-115 User Manual.

//module sdram_top (SW, KEY, CLOCK_50, LEDG, DRAM_CLK, DRAM_CKE,DRAM_ADDR, DRAM_BA, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,DRAM_WE_N, DRAM_DQ, DRAM_DQM);
module sdram_top (SW, CLOCK_50, LEDG, DRAM_CLK, DRAM_CKE,DRAM_ADDR, DRAM_BA, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,DRAM_WE_N, DRAM_DQ, DRAM_DQM);
    input[7:0]  SW;
//    input[0:0]  KEY;
    input CLOCK_50;
    output[7:0]  LEDG;
    output[12:0]  DRAM_ADDR;
    output[1:0] DRAM_BA;
    output DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK;
    output DRAM_CKE, DRAM_CS_N, DRAM_WE_N;
    output[3:0]  DRAM_DQM;
    inout[31:0]  DRAM_DQ;

// Instantiate the Nios II system module generated by the Platform Designer tool
    nios_system  NiosII  (
        .clk_clk (CLOCK_50),
//        .reset_reset_n (KEY[0]),
        .switches_export (SW),
        .leds_export (LEDG),
        .sdram_wire_addr (DRAM_ADDR),
        .sdram_wire_ba (DRAM_BA),
        .sdram_wire_cas_n (DRAM_CAS_N),
        .sdram_wire_cke (DRAM_CKE),
        .sdram_wire_cs_n (DRAM_CS_N),
        .sdram_wire_dq (DRAM_DQ),
        .sdram_wire_dqm (DRAM_DQM),
        .sdram_wire_ras_n (DRAM_RAS_N),
        .sdram_wire_we_n (DRAM_WE_N)
    );
    assignDRAM_CLK = CLOCK_50;
endmodule
