-- hw adaptation for DE1SoC Board
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY DE1SOC_COUNTER IS
GENERIC( N : INTEGER := 3 );
PORT( CLK_50 : IN STD_LOGIC
    ; KEY_RST : IN STD_LOGIC
    ; LED_COMPLETE_TICK : OUT STD_LOGIC
    ; LED_COUNT : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END DE1SOC_COUNTER;

ARCHITECTURE DE1SOC OF DE1SOC_COUNTER IS
    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';
    SIGNAL COMPLETE_TICK : STD_LOGIC := '0';
    SIGNAL COUNT : STD_LOGIC_VECTOR(N-1 DOWNTO 0) := (OTHERS => '0');

BEGIN

    COUNTER_UNIT : ENTITY
        GENERIC MAP (N => N);
        PORT MAP (CLK => CLK, RST => RST, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

    -- IN
    CLK <= CLK_50;
    RST <= NOT KEY_RST;

    -- OUT
    LED_COMPLETE_TICK <= COMPLETE_TICK;
    LED_COUNT <= COUNT;
END DE1SOC;
