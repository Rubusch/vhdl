--
-- DECODER FOR ALU
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DECODER_ENT IS
PORT( F : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; SEL : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END ENTITY DECODER_ENT;

ARCHITECTURE DECODER_ARCH OF DECODER_ENT IS
BEGIN
    SEL(0) <= F(0) AND F(1);
    SEL(1) <= F(0) AND NOT F(1);
    SEL(2) <= NOT F(0) AND F(1);
    SEL(3) <= NOT F(0) AND NOT F(1);
END ARCHITECTURE DECODER_ARCH;
