-- tb: decoder
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_DECODER IS
END TB_DECODER;

ARCHITECTURE TB OF TB_DECODER IS
    SIGNAL A : STD_LOGIC := '0';
    SIGNAL B : STD_LOGIC := '0';
    SIGNAL C : STD_LOGIC := '0';
    SIGNAL D : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    SIGNAL D_EXPECT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
    FILE INPUT_BUF : TEXT;
    FILE OUTPUT_BUF : TEXT;

BEGIN

    DECODER_UNIT : ENTITY WORK.DECODER
        PORT MAP (A => A, B => B, C => C, D => D);

    PROCESS
        VARIABLE READ_COL_FROM_INPUT_BUF : LINE;
        VARIABLE WRITE_COL_TO_OUTPUT_BUF : LINE;
        VARIABLE SEPARATOR : CHARACTER;
        VARIABLE GOOD_NUM : BOOLEAN;
        VARIABLE INPUT_A : STD_LOGIC;
        VARIABLE INPUT_B : STD_LOGIC;
        VARIABLE INPUT_C : STD_LOGIC;
        VARIABLE INPUT_D : STD_LOGIC_VECTOR(7 DOWNTO 0);
    BEGIN
        FILE_OPEN(INPUT_BUF, "../../tb_input.csv", READ_MODE);
        FILE_OPEN(OUTPUT_BUF, "../../tb_results.csv", WRITE_MODE);

        WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("A,B,C,D,D_EXPECT,TESTED"));
        WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        WHILE NOT ENDFILE(INPUT_BUF) LOOP
            READLINE(INPUT_BUF, READ_COL_FROM_INPUT_BUF);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_A, GOOD_NUM);
            NEXT WHEN NOT GOOD_NUM; --skip header

            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_B, GOOD_NUM);
            ASSERT GOOD_NUM
                REPORT("FAILURE! assignment of INPUT_B failed");
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_B);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_C);
            READ(READ_COL_FROM_INPUT_BUF, SEPARATOR);
            READ(READ_COL_FROM_INPUT_BUF, INPUT_D);

            A <= INPUT_A;
            B <= INPUT_B;
            C <= INPUT_C;
            D_EXPECT <= INPUT_D;

            WAIT FOR 20 NS;

            WRITE(WRITE_COL_TO_OUTPUT_BUF, A);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, B);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, C);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, D);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            WRITE(WRITE_COL_TO_OUTPUT_BUF, D_EXPECT);
            WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'(","));
            IF (D = D_EXPECT) THEN
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("OK"));
            ELSE
                WRITE(WRITE_COL_TO_OUTPUT_BUF, STRING'("FAIL"));
            END IF;
            WRITELINE(OUTPUT_BUF, WRITE_COL_TO_OUTPUT_BUF);

        END LOOP;
        FILE_CLOSE(INPUT_BUF);
        FILE_CLOSE(OUTPUT_BUF);
        WAIT;
    END PROCESS;
END TB;
