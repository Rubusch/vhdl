-- de1soc: hw adator for clocked shift register
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DE1SOC_SHIFTREGISTER IS
GENERIC( NBITS : INTEGER := 8);
PORT( CLK50 : IN STD_LOGIC
    ; KEY_RST : IN STD_LOGIC
    ; SW_DATA : IN STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
    ; SW_CTRL : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; LED_Q_REG : OUT STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
);
END DE1SOC_SHIFTREGISTER;

ARCHITECTURE DE1SOC OF DE1SOC_SHIFTREGISTER IS
    SIGNAL PULSE : STD_LOGIC := '0';
    SIGNAL CLK : STD_LOGIC := '0';
    SIGNAL RST : STD_LOGIC := '0';

BEGIN

    PULSE <= CLK;
    RST <= NOT KEY_RST;

    CLOCKSCALER_UNIT : ENTITY WORK.CLOCKSCALER
        GENERIC MAP (MODULO => 50000000, NBITS => 26)
        PORT MAP (CLK => CLK50, RST => RST, PULSE => PULSE);

    SHIFTREGISTER_UNIT : ENTITY WORK.SHIFTREGISTER
        GENERIC MAP (NBITS => NBITS)
        PORT MAP (CLK => CLK, RST => RST, DATA => SW_DATA, CTRL => SW_CTRL, Q_REG => LED_Q_REG);
END DE1SOC;
