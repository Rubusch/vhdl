-- de1soc: hw adapter for single port ram
--
-- author: Lothar Rubusch
-- original from: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_SINGLEPORTRAM IS
GENERIC( ADDR_WIDTH : INTEGER := 2
    ; DATA_WIDTH : INTEGER := 3
);
PORT( CLK50 : IN STD_LOGIC
    ; SW_WE : IN STD_LOGIC
    ; SW_ADDR : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; SW_DIN : IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
    ; LED_DOUT : OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
);
END DE1SOC_SINGLEPORTRAM;

ARCHITECTURE DE1SOC OF DE1SOC_SINGLEPORTRAM IS

BEGIN

    SINGLEPORTRAM_UNIT : ENTITY WORK.SINGLEPORTRAM
        PORT MAP (CLK => CLK50, WE => SW_WE, ADDR => SW_ADDR, DIN => SW_DIN, DOUT => LED_DOUT);

END DE1SOC;
