-- dual port ram
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DUALPORTRAM IS
GENERIC( ADDR_WIDTH : INTEGER := 2
    ; DATA_WIDTH : INTEGER := 3
);
PORT( CLK : IN STD_LOGIC
    ; WE : IN STD_LOGIC
    ; ADDR_WR : IN STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0)
    ; ADDR_RD : IN STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0)
    ; DIN : IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
    ; DOUT : OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
);
END DUALPORTRAM;

ARCHITECTURE DUALPORTRAM_ARCH OF DUALPORTRAM IS
    TYPE RAM_TYPE IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
    SIGNAL RAM_DUAL_PORT : RAM_TYPE;

BEGIN

    PROCESS(CLK)
    BEGIN
        IF (CLK'EVENT AND CLK = '1') THEN
            IF (WE = '1') THEN -- write data to ADDR_WR
                -- convert ADDR_WR to INTEGER from STD_LOGIC_VECTOR
                RAM_DUAL_PORT(TO_INTEGER(UNSIGNED(ADDR_WR))) <= DIN;
            ELSE
                NULL;
            END IF;
        ELSE
            NULL;
        END IF;
    END PROCESS;

    -- get address for reading data from ADDR_RD
    -- convert ADDR_RD type to INTEGER from STD_LOGIC_VECTOR
    DOUT <= RAM_DUAL_PORT(TO_INTEGER(UNSIGNED(ADDR_RD)));
END DUALPORTRAM_ARCH;
