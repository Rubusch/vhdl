--
-- A SIMPLE D-FLIPFLOP DEMO
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFLIPFLOP_ENT IS
PORT( CLK : IN STD_LOGIC
    ; RST : IN STD_LOGIC
	; D : IN STD_LOGIC
	; Q : OUT STD_LOGIC := '0'
	; QBAR : OUT STD_LOGIC := '1'
);
END ENTITY DFLIPFLOP_ENT;

ARCHITECTURE DFLIPFLOP_ARCH OF DFLIPFLOP_ENT IS

BEGIN

    P1 : PROCESS(CLK, RST)
    BEGIN
        IF RST = '0' THEN
            Q <= '0';
            QBAR <= '0';
        ELSIF (CLK'EVENT AND CLK = '1' AND RST = '1') THEN
            Q <= D;
            QBAR <= NOT D;
        END IF;
    END PROCESS;

END ARCHITECTURE DFLIPFLOP_ARCH;
