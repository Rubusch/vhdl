-- hw adaptation for DE1SoC Board: d-flipflop
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_DFLIPFLOP IS
PORT( CLK50 : IN STD_LOGIC
    ; KEY : IN STD_LOGIC
    ; SW_ENA : IN STD_LOGIC
    ; SW_D : IN STD_LOGIC
    ; LED : OUT STD_LOGIC
);
END DE1SOC_DFLIPFLOP;

ARCHITECTURE DE1SOC OF DE1SOC_DFLIPFLOP IS
    SIGNAL CLK, RST, ENA, D, Q : STD_LOGIC;

BEGIN

    DFLIPFLOP_UNIT : ENTITY WORK.DFLIPFLOP
        PORT MAP (CLK => CLK, RST => RST, ENA => ENA, D => D, Q => Q);

    -- IN
    CLK <= CLK50;
    RST <= NOT KEY;
    ENA <= SW_ENA;
    D <= SW_D;

    -- OUT
    LED <= Q;
END DE1SOC;
