-- hw adaptation for DE1SoC Board: mod-n-counter
-- (visual verification)
--
-- Author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_MODCOUNTER IS
GENERIC( NBITS : INTEGER := 2
    ; MAX_NUM : INTEGER := 4
);
PORT( CLK50 : IN STD_LOGIC
    ; KEY : IN STD_LOGIC
    ; LED : OUT STD_LOGIC
    ; LEDR : OUT STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)
);
END DE1SOC_MODCOUNTER;

ARCHITECTURE HW OF DE1SOC_MODCOUNTER IS
    SIGNAL RST : STD_LOGIC;
    SIGNAL COMPLETE_TICK : STD_LOGIC;
    SIGNAL COUNT : STD_LOGIC_VECTOR(NBITS-1 DOWNTO 0)

BEGIN

    MODCOUNTER_UNIT : ENTITY WORK.MODCOUNTER
        GENERIC MAP (NBITS => NBITS, MAX_NUM => MAX_NUM)
        PORT MAP (CLK => CLK, RST => RST, COMPLETE_TICK => COMPLETE_TICK, COUNT => COUNT);

    -- IN
    CLK <= CLK50;
    RST <= NOT KEY;

    -- OUT
    LED <= COMPLETE_TICK;
    LEDR <= COUNT;
END HW;
