--
-- FINITE STATE MACHINE (FSM) EXAMPLE
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FSM_ENT IS
PORT( RST : IN STD_LOGIC
    ; CLK : IN STD_LOGIC
    ; KEY : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; LED : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
);
END ENTITY FSM_ENT;

ARCHITECTURE FSM_ARCH OF FSM_ENT IS

BEGIN



END ARCHITECTURE FSM_ARCH;
