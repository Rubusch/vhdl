LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_NUMERIC.ALL;

ENTITY SEVENSEG_ENT IS
PORT( DATA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEG : OUT STD_LOGIC_VECTOR(13 DOWNTO 0));
END ENTITY SEVENSEG_ENT;

ARCHITECTURE SEVENSEG_ARCH OF SEVENSEG_ENT IS
BEGIN
	WITH DATA SELECT
		SEG <= "00000001111110" WHEN "0000",  -- 00
			   "00000000110000" WHEN "0001",  -- 01
			   "00000001101101" WHEN "0001",  -- 02
			   "00000001111001" WHEN "0001",  -- 03
			   "00000000110011" WHEN "0001",  -- 04
			   "00000001011011" WHEN "0001",  -- 05
--			   "0000000" WHEN "0001",  -- 06
--			   "0000000" WHEN "0001",  -- 07
--			   "0000000" WHEN "0001",  -- 08
--			   "0000000" WHEN "0001",  -- 09
--			   "01100001111110" WHEN "0001",  -- 10
--			   "" WHEN "0001",  -- 11
--			   "" WHEN "0001",  -- 12
--			   "" WHEN "0001",  -- 13
--			   "" WHEN "0001",  -- 14
--			   "" WHEN "0001",  -- 15
			   "11111101111110" WHEN OTHERS;
END ARCHITECTURE SEVENSEG_ARCH;