// nios2_hello_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2_hello_tb (
	);

	wire    nios2_hello_inst_clk_bfm_clk_clk; // nios2_hello_inst_clk_bfm:clk -> nios2_hello_inst:clk_clk

	nios2_hello nios2_hello_inst (
		.clk_clk (nios2_hello_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios2_hello_inst_clk_bfm (
		.clk (nios2_hello_inst_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
