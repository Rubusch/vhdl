-- testbench: andnand
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY TB_ANDNAND IS
PORT(
-- TODO
);
END TB_ANDNAND;

ARCHITECTURE TB OF TB_ANDNAND IS
    -- TODO
BEGIN
    -- TODO
END TB;

