--
-- LOGICAL UNIT FOR ALU
--

-- TODO