-- hw adapter: half-adder
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY DE1SOC_HALFADDER IS
PORT( SW_A : IN STD_LOGIC
    ; SW_B : IN STD_LOGIC
    ; LED_CARRY : OUT STD_LOGIC
    ; LED_SUM : OUT STD_LOGIC
);
END DE1SOC_HALFADDER;

ARCHITECTURE DE1SOC OF DE1SOC_HALFADDER IS
    SIGNAL A : STD_LOGIC := '0';
    SIGNAL B : STD_LOGIC := '0';
    SIGNAL CARRY : STD_LOGIC := '0';
    SIGNAL SUM : STD_LOGIC := '0';

BEGIN

    HALFADDER_UNIT : ENTITY WORK.HALFADDER
        PORT MAP (A => A, B => B, CARRY => CARRY, SUM => SUM);

    -- IN
    A <= SW_A;
    B <= SW_B;

    -- OUT
    LED_CARRY <= CARRY;
    LED_SUM <= SUM;
END DE1SOC;
