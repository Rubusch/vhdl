-- mod counter as state machine
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FSMCOUNTER IS
GENERIC( MODULO : NATURAL := 6
    ; NBITS : NATURAL := 4
);
PORT( CLK : IN STD_LOGIC
    ; RST : IN STD_LOGIC
    ; OUT_MOORE : OUT STD_LOGIC_VECTOR(NBITES-1 DOWNTO 0);
);
END FSMCOUNTER;

ARCHITECTURE FSM OF FSMCOUNTER IS
    TYPE STATETYPE_MOORE (START_MOORE, COUNT_MOORE);
    SIGNAL STATE_MOORE_REG, STATE_MOORE_NEXT : STATETYPE_MOORE;
    SIGNAL COUNT_MOORE_REG, COUNT_MOORE_NEXT : UNSIGNED(NBITS-1 DOWNTO 0);

BEGIN

-- TODO
END FSM
