-- hw adaptation: de1soc for alu
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_ALU IS
PORT( SW_INVA : IN STD_LOGIC
    ; SW_A : IN STD_LOGIC
    ; SW_ENA : IN STD_LOGIC
    ; SW_B : IN STD_LOGIC
    ; SW_ENB : IN STD_LOGIC
    ; SW_F : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
    ; SW_CARRY_IN : IN STD_LOGIC
    ; LED_CARRY_OUT : OUT STD_LOGIC
    ; LED_OUTPUT : OUT STD_LOGIC
);
END DE1SOC_ALU;

ARCHITECTURE DE1SOC OF DE1SOC_ALU IS
    SIGNAL INVA : STD_LOGIC := '0';
    SIGNAL A : STD_LOGIC := '0';
    SIGNAL ENA : STD_LOGIC := '0';
    SIGNAL B : STD_LOGIC := '0';
    SIGNAL ENB : STD_LOGIC := '0';
    SIGNAL F : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL CARRY_IN : STD_LOGIC := '0';
    SIGNAL CARRY_OUT : STD_LOGIC := '0';
    SIGNAL OUTPUT := STD_LOGIC := '0';

BEGIN

    ALU_UNIT : ENTITY WORK.ALU
        PORT MAP (INVA => INVA, A => A, ENA => ENA, B => B, ENB => ENB, F => F, CARRY_IN => CARRY_IN, CARRY_OUT => CARRY_OUT, OUTPUT => OUTPUT);

    -- IN
    INVA <= SW_INVA;
    A <= SW_A;
    ENA <= SW_ENA;
    B <= SW_B;
    ENB <= SW_ENB;
    F <= SW_F;
    CARRY_IN <= SW_CARRY_IN;

    -- OUT
    LED_CARRY_OUT <= CARRY_OUT;
    LED_OUTPUT <= OUTPUT;
END DE1SOC;
