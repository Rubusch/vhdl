-- testscreen: display four squares of different color on the screen
--
-- author: Lothar Rubusch
-- original from: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_TESTSCREEN IS
GENERIC();
PORT();
END DE1SOC_TESTSCREEN;

ARCHITECTURE DE1SOC OF DE1SOC_TESTSCREEN IS

BEGIN

END DE1SOC;
