-- dual port ram
--
-- author: Lothar Rubusch
-- based on: https://vhdlguide.readthedocs.io/en/latest by Meher Krishna Patel

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DUALPORTRAM IS
GENERIC();
PORT();
END DUALPORTRAM;

ARCHITECTURE DUALPORTRAM_ARCH OF DUALPORTRAM IS

BEGIN

END DUALPORTRAM_ARCH;
