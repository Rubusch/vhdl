-- HALFADDER.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HALFADDER IS
PORT( A, B : IN STD_LOGIC
    ; SUM, CARRY : OUT STD_LOGIC
    );
END HALFADDER;

ARCHITECTURE HALFADDER_ARCH OF HALFADDER IS
BEGIN
    SUM <= A XOR B;
    CARRY <= A AND B;
END HALFADDER_ARCH;
