-- hw adapter for de1soc
--
-- author: Lothar Rubusch

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE1SOC_MULTIPLEXER IS
GENERIC(NBIT : INTEGER := 4);
PORT( SW_A : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0)
    ; SW_B : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0)
    ; SW_SEL : IN STD_LOGIC
    ; LED_C : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0)
);
END DE1SOC_MULTIPLEXER;

ARCHITECTURE DE1SOC OF DE1SOC_MULTIPLEXER IS
    SIGNAL A : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL B : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL SEL : STD_LOGIC := '0';
    SIGNAL C : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0) := (OTHERS => '0');

BEGIN

    MULTIPLEXER_UNIT : ENTITY WORK.QUADMUX
        GENERIC MAP (NBIT => NBIT)
        PORT MAP (A => A, B => B, SEL => SEL, C => C);

    -- IN
    A <= SW_A;
    B <= SW_B;
    SEL <= SW_SEL;

    -- OUT
    LED_C <= C;
END DE1SOC;
